magic
tech sky130A
magscale 1 2
timestamp 1713353161
<< error_s >>
rect 20758 7946 20816 7952
rect 20950 7946 21008 7952
rect 21142 7946 21200 7952
rect 21334 7946 21392 7952
rect 21526 7946 21584 7952
rect 20758 7912 20770 7946
rect 20950 7912 20962 7946
rect 21142 7912 21154 7946
rect 21334 7912 21346 7946
rect 21526 7912 21538 7946
rect 20758 7906 20816 7912
rect 20950 7906 21008 7912
rect 21142 7906 21200 7912
rect 21334 7906 21392 7912
rect 21526 7906 21584 7912
rect 20662 6818 20720 6824
rect 20854 6818 20912 6824
rect 21046 6818 21104 6824
rect 21238 6818 21296 6824
rect 21430 6818 21488 6824
rect 20662 6784 20674 6818
rect 20854 6784 20866 6818
rect 21046 6784 21058 6818
rect 21238 6784 21250 6818
rect 21430 6784 21442 6818
rect 20662 6778 20720 6784
rect 20854 6778 20912 6784
rect 21046 6778 21104 6784
rect 21238 6778 21296 6784
rect 21430 6778 21488 6784
rect 20650 6178 20708 6184
rect 20842 6178 20900 6184
rect 21034 6178 21092 6184
rect 21226 6178 21284 6184
rect 21418 6178 21476 6184
rect 20650 6144 20662 6178
rect 20842 6144 20854 6178
rect 21034 6144 21046 6178
rect 21226 6144 21238 6178
rect 21418 6144 21430 6178
rect 20650 6138 20708 6144
rect 20842 6138 20900 6144
rect 21034 6138 21092 6144
rect 21226 6138 21284 6144
rect 21418 6138 21476 6144
rect 20746 5268 20804 5274
rect 20938 5268 20996 5274
rect 21130 5268 21188 5274
rect 21322 5268 21380 5274
rect 21514 5268 21572 5274
rect 20746 5234 20758 5268
rect 20938 5234 20950 5268
rect 21130 5234 21142 5268
rect 21322 5234 21334 5268
rect 21514 5234 21526 5268
rect 20746 5228 20804 5234
rect 20938 5228 20996 5234
rect 21130 5228 21188 5234
rect 21322 5228 21380 5234
rect 21514 5228 21572 5234
rect 20746 5160 20804 5166
rect 20938 5160 20996 5166
rect 21130 5160 21188 5166
rect 21322 5160 21380 5166
rect 21514 5160 21572 5166
rect 20746 5126 20758 5160
rect 20938 5126 20950 5160
rect 21130 5126 21142 5160
rect 21322 5126 21334 5160
rect 21514 5126 21526 5160
rect 20746 5120 20804 5126
rect 20938 5120 20996 5126
rect 21130 5120 21188 5126
rect 21322 5120 21380 5126
rect 21514 5120 21572 5126
rect 20650 4250 20708 4256
rect 20842 4250 20900 4256
rect 21034 4250 21092 4256
rect 21226 4250 21284 4256
rect 21418 4250 21476 4256
rect 20650 4216 20662 4250
rect 20842 4216 20854 4250
rect 21034 4216 21046 4250
rect 21226 4216 21238 4250
rect 21418 4216 21430 4250
rect 20650 4210 20708 4216
rect 20842 4210 20900 4216
rect 21034 4210 21092 4216
rect 21226 4210 21284 4216
rect 21418 4210 21476 4216
rect 7987 3874 8045 3880
rect 8105 3874 8163 3880
rect 8223 3874 8281 3880
rect 8341 3874 8399 3880
rect 8459 3874 8517 3880
rect 8577 3874 8635 3880
rect 8695 3874 8753 3880
rect 8813 3874 8871 3880
rect 8931 3874 8989 3880
rect 9049 3874 9107 3880
rect 9167 3874 9225 3880
rect 9285 3874 9343 3880
rect 9403 3874 9461 3880
rect 9521 3874 9579 3880
rect 9639 3874 9697 3880
rect 9757 3874 9815 3880
rect 9875 3874 9933 3880
rect 9993 3874 10051 3880
rect 10111 3874 10169 3880
rect 10229 3874 10287 3880
rect 7987 3840 7999 3874
rect 8105 3840 8117 3874
rect 8223 3840 8235 3874
rect 8341 3840 8353 3874
rect 8459 3840 8471 3874
rect 8577 3840 8589 3874
rect 8695 3840 8707 3874
rect 8813 3840 8825 3874
rect 8931 3840 8943 3874
rect 9049 3840 9061 3874
rect 9167 3840 9179 3874
rect 9285 3840 9297 3874
rect 9403 3840 9415 3874
rect 9521 3840 9533 3874
rect 9639 3840 9651 3874
rect 9757 3840 9769 3874
rect 9875 3840 9887 3874
rect 9993 3840 10005 3874
rect 10111 3840 10123 3874
rect 10229 3840 10241 3874
rect 7987 3834 8045 3840
rect 8105 3834 8163 3840
rect 8223 3834 8281 3840
rect 8341 3834 8399 3840
rect 8459 3834 8517 3840
rect 8577 3834 8635 3840
rect 8695 3834 8753 3840
rect 8813 3834 8871 3840
rect 8931 3834 8989 3840
rect 9049 3834 9107 3840
rect 9167 3834 9225 3840
rect 9285 3834 9343 3840
rect 9403 3834 9461 3840
rect 9521 3834 9579 3840
rect 9639 3834 9697 3840
rect 9757 3834 9815 3840
rect 9875 3834 9933 3840
rect 9993 3834 10051 3840
rect 10111 3834 10169 3840
rect 10229 3834 10287 3840
rect 7987 3364 8045 3370
rect 8105 3364 8163 3370
rect 8223 3364 8281 3370
rect 8341 3364 8399 3370
rect 8459 3364 8517 3370
rect 8577 3364 8635 3370
rect 8695 3364 8753 3370
rect 8813 3364 8871 3370
rect 8931 3364 8989 3370
rect 9049 3364 9107 3370
rect 9167 3364 9225 3370
rect 9285 3364 9343 3370
rect 9403 3364 9461 3370
rect 9521 3364 9579 3370
rect 9639 3364 9697 3370
rect 9757 3364 9815 3370
rect 9875 3364 9933 3370
rect 9993 3364 10051 3370
rect 10111 3364 10169 3370
rect 10229 3364 10287 3370
rect 7987 3330 7999 3364
rect 8105 3330 8117 3364
rect 8223 3330 8235 3364
rect 8341 3330 8353 3364
rect 8459 3330 8471 3364
rect 8577 3330 8589 3364
rect 8695 3330 8707 3364
rect 8813 3330 8825 3364
rect 8931 3330 8943 3364
rect 9049 3330 9061 3364
rect 9167 3330 9179 3364
rect 9285 3330 9297 3364
rect 9403 3330 9415 3364
rect 9521 3330 9533 3364
rect 9639 3330 9651 3364
rect 9757 3330 9769 3364
rect 9875 3330 9887 3364
rect 9993 3330 10005 3364
rect 10111 3330 10123 3364
rect 10229 3330 10241 3364
rect 7987 3324 8045 3330
rect 8105 3324 8163 3330
rect 8223 3324 8281 3330
rect 8341 3324 8399 3330
rect 8459 3324 8517 3330
rect 8577 3324 8635 3330
rect 8695 3324 8753 3330
rect 8813 3324 8871 3330
rect 8931 3324 8989 3330
rect 9049 3324 9107 3330
rect 9167 3324 9225 3330
rect 9285 3324 9343 3330
rect 9403 3324 9461 3330
rect 9521 3324 9579 3330
rect 9639 3324 9697 3330
rect 9757 3324 9815 3330
rect 9875 3324 9933 3330
rect 9993 3324 10051 3330
rect 10111 3324 10169 3330
rect 10229 3324 10287 3330
<< pwell >>
rect 1872 7070 1982 7542
rect 2684 7472 2800 7944
rect 5588 7716 7106 7774
rect 5588 7398 7106 7456
rect 5588 7300 7106 7358
rect 5588 6982 7106 7040
rect 5588 6884 7106 6942
rect 5588 6566 7106 6624
rect 5588 6462 7106 6520
rect 5588 6146 7106 6204
rect 5594 6046 7112 6104
rect 5588 5730 7106 5788
rect 2564 2372 2632 2528
rect 3484 2372 3552 2528
rect 4398 2372 4466 2528
rect 5314 2372 5382 2528
<< viali >>
rect 4352 9918 4562 9988
rect 6330 9916 6522 9984
rect 8164 9936 8432 10006
rect 12314 9934 12618 10008
rect 14222 9936 14510 10006
rect 18376 9932 18668 10008
rect 20274 9878 20448 9954
rect 21366 9880 21528 9956
rect 1078 4942 1242 4998
rect 1472 4942 1636 4998
rect 1866 4942 2030 4998
rect 2258 4942 2428 5000
rect 2670 4942 2834 5000
rect 3062 4942 3224 5000
rect 1068 3292 1142 3556
rect 2038 2042 2246 2134
rect 4814 2046 5046 2134
rect 7516 2052 7754 2138
rect 10260 2052 10500 2136
rect 12758 2052 12986 2138
rect 15548 2054 15776 2136
rect 17912 2060 18164 2136
rect 20726 2056 20964 2136
<< metal1 >>
rect 30 10348 22606 10794
rect 546 10136 752 10348
rect 546 9924 752 9930
rect 4312 9988 4604 10348
rect 4312 9918 4352 9988
rect 4562 9918 4604 9988
rect 4312 9908 4604 9918
rect 6276 9984 6568 10348
rect 6276 9916 6330 9984
rect 6522 9916 6568 9984
rect 8088 10006 8492 10348
rect 8088 9936 8164 10006
rect 8432 9936 8492 10006
rect 8088 9922 8492 9936
rect 12264 10008 12668 10348
rect 12264 9934 12314 10008
rect 12618 9934 12668 10008
rect 12264 9920 12668 9934
rect 14158 10006 14562 10348
rect 14158 9936 14222 10006
rect 14510 9936 14562 10006
rect 14158 9924 14562 9936
rect 18324 10008 18728 10348
rect 18324 9932 18376 10008
rect 18668 9932 18728 10008
rect 18324 9922 18728 9932
rect 20240 9954 20478 10348
rect 6276 9906 6568 9916
rect 20240 9878 20274 9954
rect 20448 9878 20478 9954
rect 20240 9870 20478 9878
rect 21332 9956 21570 10348
rect 21332 9880 21366 9956
rect 21528 9880 21570 9956
rect 21332 9866 21570 9880
rect 102 8284 3830 8484
rect 3630 8096 3830 8284
rect 2293 7542 2403 7941
rect 1128 7436 1610 7536
rect 540 6937 546 7143
rect 752 6937 758 7143
rect 1128 7074 1222 7436
rect 1510 7080 1610 7436
rect 1872 7432 2403 7542
rect 2684 7828 3202 7944
rect 2684 7472 2800 7828
rect 3086 7450 3202 7828
rect 3658 7774 3803 8096
rect 3658 7716 5226 7774
rect 5588 7716 7106 7774
rect 3658 7714 3803 7716
rect 3708 7456 3766 7714
rect 7045 7456 7103 7716
rect 1872 7070 1982 7432
rect 3708 7398 5226 7456
rect 5588 7398 7106 7456
rect 3708 7358 3766 7398
rect 7045 7358 7103 7398
rect 3708 7300 5226 7358
rect 5588 7300 7106 7358
rect 3708 7040 3766 7300
rect 7045 7040 7103 7300
rect 3708 6982 5226 7040
rect 5588 6982 7106 7040
rect 3708 6942 3766 6982
rect 7045 6942 7103 6982
rect 546 5338 752 6937
rect 3708 6884 5226 6942
rect 5588 6884 7106 6942
rect 3708 6624 3766 6884
rect 7045 6624 7103 6884
rect 3708 6566 5226 6624
rect 5588 6566 7106 6624
rect 3708 6520 3766 6566
rect 7045 6520 7103 6566
rect 3708 6462 5226 6520
rect 5588 6462 7106 6520
rect 3708 6204 3766 6462
rect 7045 6204 7103 6462
rect 22378 6402 22578 6602
rect 3708 6146 5226 6204
rect 5588 6146 7106 6204
rect 3708 6104 3766 6146
rect 7045 6104 7103 6146
rect 3708 6046 5226 6104
rect 5594 6046 7112 6104
rect 3708 5788 3766 6046
rect 7045 5788 7103 6046
rect 3708 5730 5226 5788
rect 5588 5730 7106 5788
rect 7045 5652 7103 5730
rect 1110 5338 1218 5538
rect 546 5132 1218 5338
rect 1502 5172 1606 5528
rect 1878 5172 1982 5524
rect 1502 5068 1982 5172
rect 2290 5178 2404 5528
rect 2689 5178 2803 5549
rect 7025 5543 7124 5652
rect 2290 5064 2803 5178
rect 3088 5174 3188 5536
rect 6989 5179 7159 5543
rect 3084 5168 3520 5174
rect 3084 5078 3636 5168
rect 3088 5075 3188 5078
rect 814 5000 3242 5014
rect 814 4998 2258 5000
rect 814 4942 1078 4998
rect 1242 4942 1472 4998
rect 1636 4942 1866 4998
rect 2030 4942 2258 4998
rect 2428 4942 2670 5000
rect 2834 4942 3062 5000
rect 3224 4942 3242 5000
rect 814 4930 3242 4942
rect 98 4358 298 4386
rect 475 4363 645 4369
rect 98 4199 475 4358
rect 98 4186 298 4199
rect 475 4187 645 4193
rect 814 3582 898 4930
rect 3428 4072 3636 5078
rect 6989 5003 7159 5009
rect 22380 4698 22580 4898
rect 1533 4002 1682 4008
rect 3428 4002 6574 4072
rect 1682 3864 6574 4002
rect 1682 3853 3678 3864
rect 1533 3847 1682 3853
rect 1218 3627 6304 3630
rect 6495 3627 6569 3864
rect 49 3556 1148 3582
rect 1218 3556 6569 3627
rect 49 3292 1068 3556
rect 1142 3292 1148 3556
rect 6255 3553 6569 3556
rect 1190 3460 1200 3522
rect 1256 3460 1266 3522
rect 2106 3460 2116 3522
rect 2172 3460 2182 3522
rect 3022 3460 3032 3522
rect 3088 3460 3098 3522
rect 3938 3460 3948 3522
rect 4004 3460 4014 3522
rect 4852 3456 4862 3518
rect 4918 3456 4928 3518
rect 5768 3458 5778 3520
rect 5834 3458 5844 3520
rect 1642 3318 1652 3374
rect 1722 3318 1732 3374
rect 2558 3318 2568 3374
rect 2638 3318 2648 3374
rect 3472 3320 3482 3376
rect 3552 3320 3562 3376
rect 4390 3318 4400 3374
rect 4470 3318 4480 3374
rect 5306 3318 5316 3374
rect 5386 3318 5396 3374
rect 49 3272 1148 3292
rect 6495 3282 6569 3553
rect 49 1528 359 3272
rect 575 3270 768 3272
rect 1222 3208 6569 3282
rect 746 2923 873 2929
rect 746 2664 873 2796
rect 6131 2789 6137 2851
rect 6199 2789 6205 2851
rect 780 2546 838 2664
rect 780 2545 5800 2546
rect 778 2488 5800 2545
rect 778 2230 828 2488
rect 1652 2372 1720 2488
rect 2564 2372 2632 2488
rect 3484 2372 3552 2488
rect 4398 2372 4466 2488
rect 5314 2372 5382 2488
rect 1180 2262 1190 2318
rect 1260 2262 1270 2318
rect 2098 2264 2108 2320
rect 2178 2264 2188 2320
rect 3012 2264 3022 2320
rect 3092 2264 3102 2320
rect 3930 2264 3940 2320
rect 4010 2264 4020 2320
rect 4844 2264 4854 2320
rect 4924 2264 4934 2320
rect 5764 2264 5774 2320
rect 5844 2264 5854 2320
rect 778 2180 5798 2230
rect 1972 2134 2310 2148
rect 1972 2042 2038 2134
rect 2246 2042 2310 2134
rect 575 1528 830 1530
rect 1972 1528 2310 2042
rect 4762 2134 5098 2148
rect 4762 2046 4814 2134
rect 5046 2046 5098 2134
rect 4762 1528 5098 2046
rect 6137 1528 6199 2789
rect 7462 2138 7800 2150
rect 7462 2052 7516 2138
rect 7754 2052 7800 2138
rect 7462 1528 7800 2052
rect 10206 2136 10546 2148
rect 10206 2052 10260 2136
rect 10500 2052 10546 2136
rect 10206 1528 10546 2052
rect 12692 2138 13036 2150
rect 12692 2052 12758 2138
rect 12986 2052 13036 2138
rect 12692 1528 13036 2052
rect 15488 2136 15834 2148
rect 15488 2054 15548 2136
rect 15776 2054 15834 2136
rect 15488 1528 15834 2054
rect 17864 2136 18210 2148
rect 17864 2060 17912 2136
rect 18164 2060 18210 2136
rect 17864 2052 18210 2060
rect 20676 2136 21024 2148
rect 20676 2056 20726 2136
rect 20964 2056 21024 2136
rect 17864 1528 18212 2052
rect 20676 1528 21024 2056
rect 10 1494 22586 1528
rect 10 1404 1000 1494
rect 1240 1404 22586 1494
rect 10 1082 22586 1404
rect 17864 1078 18212 1082
<< via1 >>
rect 546 9930 752 10136
rect 546 6937 752 7143
rect 475 4193 645 4363
rect 6989 5009 7159 5179
rect 1533 3853 1682 4002
rect 1200 3460 1256 3522
rect 2116 3460 2172 3522
rect 3032 3460 3088 3522
rect 3948 3460 4004 3522
rect 4862 3456 4918 3518
rect 5778 3458 5834 3520
rect 1652 3318 1722 3374
rect 2568 3318 2638 3374
rect 3482 3320 3552 3376
rect 4400 3318 4470 3374
rect 5316 3318 5386 3374
rect 746 2796 873 2923
rect 6137 2789 6199 2851
rect 1190 2262 1260 2318
rect 2108 2264 2178 2320
rect 3022 2264 3092 2320
rect 3940 2264 4010 2320
rect 4854 2264 4924 2320
rect 5774 2264 5844 2320
rect 1000 1404 1240 1494
<< metal2 >>
rect 540 9930 546 10136
rect 752 9930 758 10136
rect 546 7143 752 9930
rect 546 6931 752 6937
rect 6983 5009 6989 5179
rect 7159 5009 7165 5179
rect 6989 4363 7159 5009
rect 469 4193 475 4363
rect 645 4193 7159 4363
rect 735 3853 1533 4002
rect 1682 3853 1688 4002
rect 746 2923 873 3853
rect 1200 3522 1256 3532
rect 2116 3522 2172 3532
rect 3032 3522 3088 3532
rect 3948 3522 4004 3532
rect 4862 3522 4918 3528
rect 5778 3522 5834 3530
rect 1182 3460 1200 3522
rect 1256 3460 2116 3522
rect 2172 3460 3032 3522
rect 3088 3460 3948 3522
rect 4004 3520 6200 3522
rect 4004 3518 5778 3520
rect 4004 3460 4862 3518
rect 1182 3458 4862 3460
rect 1200 3450 1256 3458
rect 2116 3450 2172 3458
rect 3032 3450 3088 3458
rect 3948 3450 4004 3458
rect 4918 3458 5778 3518
rect 5834 3458 6200 3520
rect 4862 3446 4918 3456
rect 5778 3448 5834 3458
rect 1652 3374 1722 3384
rect 2568 3374 2638 3384
rect 3482 3376 3552 3386
rect 1180 3318 1652 3374
rect 1722 3318 2568 3374
rect 2638 3320 3482 3374
rect 4400 3374 4470 3384
rect 5316 3374 5386 3384
rect 3552 3320 4400 3374
rect 2638 3318 4400 3320
rect 4470 3318 5316 3374
rect 5386 3318 6200 3374
rect 1180 3312 6200 3318
rect 1652 3308 1722 3312
rect 2568 3308 2638 3312
rect 3482 3310 3552 3312
rect 4400 3308 4470 3312
rect 5316 3308 5386 3312
rect 740 2796 746 2923
rect 873 2796 879 2923
rect 6137 2851 6199 3312
rect 6137 2783 6199 2789
rect 1190 2318 1260 2328
rect 912 2262 1190 2312
rect 2108 2320 2178 2330
rect 1260 2264 2108 2312
rect 3022 2320 3092 2330
rect 2178 2264 3022 2312
rect 3940 2320 4010 2330
rect 3092 2264 3940 2312
rect 4854 2320 4924 2330
rect 4010 2264 4854 2312
rect 5774 2320 5844 2330
rect 4924 2264 5774 2312
rect 5844 2264 5860 2312
rect 1260 2262 5860 2264
rect 912 2252 5860 2262
rect 912 1480 972 2252
rect 1000 1494 1240 1504
rect 912 1420 1000 1480
rect 1000 1394 1240 1404
use sky130_fd_pr__nfet_01v8_FMJ72H  XM1
timestamp 1713266475
transform 1 0 4651 0 1 6752
box -757 -1146 757 1146
use sky130_fd_pr__nfet_01v8_FMJ72H  XM2
timestamp 1713266475
transform 1 0 6159 0 1 6752
box -757 -1146 757 1146
use sky130_fd_pr__pfet_01v8_3H5TVM  XM3
timestamp 1713266475
transform 1 0 6410 0 1 9677
box -812 -319 812 319
use sky130_fd_pr__pfet_01v8_3H5TVM  XM4
timestamp 1713266475
transform 1 0 4454 0 1 9683
box -812 -319 812 319
use sky130_fd_pr__nfet_01v8_EPHDNF  XM5
timestamp 1713266475
transform 1 0 3517 0 1 3420
box -2457 -310 2457 310
use sky130_fd_pr__nfet_01v8_EPHDNF  XM6
timestamp 1713266475
transform 1 0 3517 0 1 2358
box -2457 -310 2457 310
use sky130_fd_pr__nfet_01v8_SMX62R  XM7
timestamp 1713266475
transform 1 0 9137 0 1 3602
box -1347 -410 1347 410
use sky130_fd_pr__nfet_01v8_EPHDNF  XM8
timestamp 1713266475
transform 1 0 8991 0 1 2356
box -2457 -310 2457 310
use sky130_fd_pr__pfet_01v8_P7N2DR  XM9
timestamp 1713266475
transform 1 0 10459 0 1 7343
box -2747 -2677 2747 2677
use sky130_fd_pr__pfet_01v8_P7N2DR  XM10
timestamp 1713266475
transform 1 0 16531 0 1 7343
box -2747 -2677 2747 2677
use sky130_fd_pr__nfet_01v8_EPHDNF  XM11
timestamp 1713266475
transform 1 0 14255 0 1 2358
box -2457 -310 2457 310
use sky130_fd_pr__nfet_01v8_V5FT3Q  XM12
timestamp 1713266475
transform 1 0 20546 0 1 3358
box -1312 -410 1312 410
use sky130_fd_pr__pfet_01v8_3HZ9VM  XM13
timestamp 1713266475
transform 1 0 20354 0 1 9245
box -296 -719 296 719
use sky130_fd_pr__nfet_01v8_EPHDNF  XM14
timestamp 1713266475
transform 1 0 19417 0 1 2358
box -2457 -310 2457 310
use sky130_fd_pr__nfet_01v8_GSBCLJ  XM15
timestamp 1713266475
transform 1 0 21111 0 1 5197
box -647 -1119 647 1119
use sky130_fd_pr__pfet_01v8_3HZ9VM  XM16
timestamp 1713266475
transform 1 0 21446 0 1 9243
box -296 -719 296 719
use sky130_fd_pr__pfet_01v8_BDVWJN  XM17
timestamp 1713266475
transform 1 0 21123 0 1 7365
box -647 -719 647 719
use sky130_fd_pr__res_xhigh_po_0p35_RF5GSL  XR1
timestamp 1713266475
transform 1 0 1553 0 1 6300
box -201 -1382 201 1382
use sky130_fd_pr__res_xhigh_po_0p35_RF5GSL  XR2
timestamp 1713266475
transform 1 0 1161 0 1 6300
box -201 -1382 201 1382
use sky130_fd_pr__res_xhigh_po_0p35_RF5GSL  XR3
timestamp 1713266475
transform 1 0 1947 0 1 6300
box -201 -1382 201 1382
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR4
timestamp 1713266475
transform 1 0 2345 0 1 6500
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR5
timestamp 1713266475
transform 1 0 3143 0 1 6500
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR6
timestamp 1713266475
transform 1 0 2749 0 1 6500
box -201 -1582 201 1582
<< labels >>
flabel metal1 106 1246 306 1446 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 22378 6402 22578 6602 0 FreeSans 256 0 0 0 z
port 2 nsew
flabel metal1 22380 4698 22580 4898 0 FreeSans 256 0 0 0 x
port 5 nsew
flabel metal1 98 4186 298 4386 0 FreeSans 256 0 0 0 y
port 3 nsew
flabel metal1 102 8284 302 8484 0 FreeSans 256 0 0 0 ref
port 4 nsew
flabel metal1 92 10506 292 10706 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 3428 3864 6574 4072 0 FreeSans 1600 0 0 0 G2
<< end >>
