magic
tech sky130A
magscale 1 2
timestamp 1713266475
<< nwell >>
rect -2747 -2677 2747 2677
<< pmos >>
rect -2551 1958 -2351 2458
rect -2293 1958 -2093 2458
rect -2035 1958 -1835 2458
rect -1777 1958 -1577 2458
rect -1519 1958 -1319 2458
rect -1261 1958 -1061 2458
rect -1003 1958 -803 2458
rect -745 1958 -545 2458
rect -487 1958 -287 2458
rect -229 1958 -29 2458
rect 29 1958 229 2458
rect 287 1958 487 2458
rect 545 1958 745 2458
rect 803 1958 1003 2458
rect 1061 1958 1261 2458
rect 1319 1958 1519 2458
rect 1577 1958 1777 2458
rect 1835 1958 2035 2458
rect 2093 1958 2293 2458
rect 2351 1958 2551 2458
rect -2551 1222 -2351 1722
rect -2293 1222 -2093 1722
rect -2035 1222 -1835 1722
rect -1777 1222 -1577 1722
rect -1519 1222 -1319 1722
rect -1261 1222 -1061 1722
rect -1003 1222 -803 1722
rect -745 1222 -545 1722
rect -487 1222 -287 1722
rect -229 1222 -29 1722
rect 29 1222 229 1722
rect 287 1222 487 1722
rect 545 1222 745 1722
rect 803 1222 1003 1722
rect 1061 1222 1261 1722
rect 1319 1222 1519 1722
rect 1577 1222 1777 1722
rect 1835 1222 2035 1722
rect 2093 1222 2293 1722
rect 2351 1222 2551 1722
rect -2551 486 -2351 986
rect -2293 486 -2093 986
rect -2035 486 -1835 986
rect -1777 486 -1577 986
rect -1519 486 -1319 986
rect -1261 486 -1061 986
rect -1003 486 -803 986
rect -745 486 -545 986
rect -487 486 -287 986
rect -229 486 -29 986
rect 29 486 229 986
rect 287 486 487 986
rect 545 486 745 986
rect 803 486 1003 986
rect 1061 486 1261 986
rect 1319 486 1519 986
rect 1577 486 1777 986
rect 1835 486 2035 986
rect 2093 486 2293 986
rect 2351 486 2551 986
rect -2551 -250 -2351 250
rect -2293 -250 -2093 250
rect -2035 -250 -1835 250
rect -1777 -250 -1577 250
rect -1519 -250 -1319 250
rect -1261 -250 -1061 250
rect -1003 -250 -803 250
rect -745 -250 -545 250
rect -487 -250 -287 250
rect -229 -250 -29 250
rect 29 -250 229 250
rect 287 -250 487 250
rect 545 -250 745 250
rect 803 -250 1003 250
rect 1061 -250 1261 250
rect 1319 -250 1519 250
rect 1577 -250 1777 250
rect 1835 -250 2035 250
rect 2093 -250 2293 250
rect 2351 -250 2551 250
rect -2551 -986 -2351 -486
rect -2293 -986 -2093 -486
rect -2035 -986 -1835 -486
rect -1777 -986 -1577 -486
rect -1519 -986 -1319 -486
rect -1261 -986 -1061 -486
rect -1003 -986 -803 -486
rect -745 -986 -545 -486
rect -487 -986 -287 -486
rect -229 -986 -29 -486
rect 29 -986 229 -486
rect 287 -986 487 -486
rect 545 -986 745 -486
rect 803 -986 1003 -486
rect 1061 -986 1261 -486
rect 1319 -986 1519 -486
rect 1577 -986 1777 -486
rect 1835 -986 2035 -486
rect 2093 -986 2293 -486
rect 2351 -986 2551 -486
rect -2551 -1722 -2351 -1222
rect -2293 -1722 -2093 -1222
rect -2035 -1722 -1835 -1222
rect -1777 -1722 -1577 -1222
rect -1519 -1722 -1319 -1222
rect -1261 -1722 -1061 -1222
rect -1003 -1722 -803 -1222
rect -745 -1722 -545 -1222
rect -487 -1722 -287 -1222
rect -229 -1722 -29 -1222
rect 29 -1722 229 -1222
rect 287 -1722 487 -1222
rect 545 -1722 745 -1222
rect 803 -1722 1003 -1222
rect 1061 -1722 1261 -1222
rect 1319 -1722 1519 -1222
rect 1577 -1722 1777 -1222
rect 1835 -1722 2035 -1222
rect 2093 -1722 2293 -1222
rect 2351 -1722 2551 -1222
rect -2551 -2458 -2351 -1958
rect -2293 -2458 -2093 -1958
rect -2035 -2458 -1835 -1958
rect -1777 -2458 -1577 -1958
rect -1519 -2458 -1319 -1958
rect -1261 -2458 -1061 -1958
rect -1003 -2458 -803 -1958
rect -745 -2458 -545 -1958
rect -487 -2458 -287 -1958
rect -229 -2458 -29 -1958
rect 29 -2458 229 -1958
rect 287 -2458 487 -1958
rect 545 -2458 745 -1958
rect 803 -2458 1003 -1958
rect 1061 -2458 1261 -1958
rect 1319 -2458 1519 -1958
rect 1577 -2458 1777 -1958
rect 1835 -2458 2035 -1958
rect 2093 -2458 2293 -1958
rect 2351 -2458 2551 -1958
<< pdiff >>
rect -2609 2446 -2551 2458
rect -2609 1970 -2597 2446
rect -2563 1970 -2551 2446
rect -2609 1958 -2551 1970
rect -2351 2446 -2293 2458
rect -2351 1970 -2339 2446
rect -2305 1970 -2293 2446
rect -2351 1958 -2293 1970
rect -2093 2446 -2035 2458
rect -2093 1970 -2081 2446
rect -2047 1970 -2035 2446
rect -2093 1958 -2035 1970
rect -1835 2446 -1777 2458
rect -1835 1970 -1823 2446
rect -1789 1970 -1777 2446
rect -1835 1958 -1777 1970
rect -1577 2446 -1519 2458
rect -1577 1970 -1565 2446
rect -1531 1970 -1519 2446
rect -1577 1958 -1519 1970
rect -1319 2446 -1261 2458
rect -1319 1970 -1307 2446
rect -1273 1970 -1261 2446
rect -1319 1958 -1261 1970
rect -1061 2446 -1003 2458
rect -1061 1970 -1049 2446
rect -1015 1970 -1003 2446
rect -1061 1958 -1003 1970
rect -803 2446 -745 2458
rect -803 1970 -791 2446
rect -757 1970 -745 2446
rect -803 1958 -745 1970
rect -545 2446 -487 2458
rect -545 1970 -533 2446
rect -499 1970 -487 2446
rect -545 1958 -487 1970
rect -287 2446 -229 2458
rect -287 1970 -275 2446
rect -241 1970 -229 2446
rect -287 1958 -229 1970
rect -29 2446 29 2458
rect -29 1970 -17 2446
rect 17 1970 29 2446
rect -29 1958 29 1970
rect 229 2446 287 2458
rect 229 1970 241 2446
rect 275 1970 287 2446
rect 229 1958 287 1970
rect 487 2446 545 2458
rect 487 1970 499 2446
rect 533 1970 545 2446
rect 487 1958 545 1970
rect 745 2446 803 2458
rect 745 1970 757 2446
rect 791 1970 803 2446
rect 745 1958 803 1970
rect 1003 2446 1061 2458
rect 1003 1970 1015 2446
rect 1049 1970 1061 2446
rect 1003 1958 1061 1970
rect 1261 2446 1319 2458
rect 1261 1970 1273 2446
rect 1307 1970 1319 2446
rect 1261 1958 1319 1970
rect 1519 2446 1577 2458
rect 1519 1970 1531 2446
rect 1565 1970 1577 2446
rect 1519 1958 1577 1970
rect 1777 2446 1835 2458
rect 1777 1970 1789 2446
rect 1823 1970 1835 2446
rect 1777 1958 1835 1970
rect 2035 2446 2093 2458
rect 2035 1970 2047 2446
rect 2081 1970 2093 2446
rect 2035 1958 2093 1970
rect 2293 2446 2351 2458
rect 2293 1970 2305 2446
rect 2339 1970 2351 2446
rect 2293 1958 2351 1970
rect 2551 2446 2609 2458
rect 2551 1970 2563 2446
rect 2597 1970 2609 2446
rect 2551 1958 2609 1970
rect -2609 1710 -2551 1722
rect -2609 1234 -2597 1710
rect -2563 1234 -2551 1710
rect -2609 1222 -2551 1234
rect -2351 1710 -2293 1722
rect -2351 1234 -2339 1710
rect -2305 1234 -2293 1710
rect -2351 1222 -2293 1234
rect -2093 1710 -2035 1722
rect -2093 1234 -2081 1710
rect -2047 1234 -2035 1710
rect -2093 1222 -2035 1234
rect -1835 1710 -1777 1722
rect -1835 1234 -1823 1710
rect -1789 1234 -1777 1710
rect -1835 1222 -1777 1234
rect -1577 1710 -1519 1722
rect -1577 1234 -1565 1710
rect -1531 1234 -1519 1710
rect -1577 1222 -1519 1234
rect -1319 1710 -1261 1722
rect -1319 1234 -1307 1710
rect -1273 1234 -1261 1710
rect -1319 1222 -1261 1234
rect -1061 1710 -1003 1722
rect -1061 1234 -1049 1710
rect -1015 1234 -1003 1710
rect -1061 1222 -1003 1234
rect -803 1710 -745 1722
rect -803 1234 -791 1710
rect -757 1234 -745 1710
rect -803 1222 -745 1234
rect -545 1710 -487 1722
rect -545 1234 -533 1710
rect -499 1234 -487 1710
rect -545 1222 -487 1234
rect -287 1710 -229 1722
rect -287 1234 -275 1710
rect -241 1234 -229 1710
rect -287 1222 -229 1234
rect -29 1710 29 1722
rect -29 1234 -17 1710
rect 17 1234 29 1710
rect -29 1222 29 1234
rect 229 1710 287 1722
rect 229 1234 241 1710
rect 275 1234 287 1710
rect 229 1222 287 1234
rect 487 1710 545 1722
rect 487 1234 499 1710
rect 533 1234 545 1710
rect 487 1222 545 1234
rect 745 1710 803 1722
rect 745 1234 757 1710
rect 791 1234 803 1710
rect 745 1222 803 1234
rect 1003 1710 1061 1722
rect 1003 1234 1015 1710
rect 1049 1234 1061 1710
rect 1003 1222 1061 1234
rect 1261 1710 1319 1722
rect 1261 1234 1273 1710
rect 1307 1234 1319 1710
rect 1261 1222 1319 1234
rect 1519 1710 1577 1722
rect 1519 1234 1531 1710
rect 1565 1234 1577 1710
rect 1519 1222 1577 1234
rect 1777 1710 1835 1722
rect 1777 1234 1789 1710
rect 1823 1234 1835 1710
rect 1777 1222 1835 1234
rect 2035 1710 2093 1722
rect 2035 1234 2047 1710
rect 2081 1234 2093 1710
rect 2035 1222 2093 1234
rect 2293 1710 2351 1722
rect 2293 1234 2305 1710
rect 2339 1234 2351 1710
rect 2293 1222 2351 1234
rect 2551 1710 2609 1722
rect 2551 1234 2563 1710
rect 2597 1234 2609 1710
rect 2551 1222 2609 1234
rect -2609 974 -2551 986
rect -2609 498 -2597 974
rect -2563 498 -2551 974
rect -2609 486 -2551 498
rect -2351 974 -2293 986
rect -2351 498 -2339 974
rect -2305 498 -2293 974
rect -2351 486 -2293 498
rect -2093 974 -2035 986
rect -2093 498 -2081 974
rect -2047 498 -2035 974
rect -2093 486 -2035 498
rect -1835 974 -1777 986
rect -1835 498 -1823 974
rect -1789 498 -1777 974
rect -1835 486 -1777 498
rect -1577 974 -1519 986
rect -1577 498 -1565 974
rect -1531 498 -1519 974
rect -1577 486 -1519 498
rect -1319 974 -1261 986
rect -1319 498 -1307 974
rect -1273 498 -1261 974
rect -1319 486 -1261 498
rect -1061 974 -1003 986
rect -1061 498 -1049 974
rect -1015 498 -1003 974
rect -1061 486 -1003 498
rect -803 974 -745 986
rect -803 498 -791 974
rect -757 498 -745 974
rect -803 486 -745 498
rect -545 974 -487 986
rect -545 498 -533 974
rect -499 498 -487 974
rect -545 486 -487 498
rect -287 974 -229 986
rect -287 498 -275 974
rect -241 498 -229 974
rect -287 486 -229 498
rect -29 974 29 986
rect -29 498 -17 974
rect 17 498 29 974
rect -29 486 29 498
rect 229 974 287 986
rect 229 498 241 974
rect 275 498 287 974
rect 229 486 287 498
rect 487 974 545 986
rect 487 498 499 974
rect 533 498 545 974
rect 487 486 545 498
rect 745 974 803 986
rect 745 498 757 974
rect 791 498 803 974
rect 745 486 803 498
rect 1003 974 1061 986
rect 1003 498 1015 974
rect 1049 498 1061 974
rect 1003 486 1061 498
rect 1261 974 1319 986
rect 1261 498 1273 974
rect 1307 498 1319 974
rect 1261 486 1319 498
rect 1519 974 1577 986
rect 1519 498 1531 974
rect 1565 498 1577 974
rect 1519 486 1577 498
rect 1777 974 1835 986
rect 1777 498 1789 974
rect 1823 498 1835 974
rect 1777 486 1835 498
rect 2035 974 2093 986
rect 2035 498 2047 974
rect 2081 498 2093 974
rect 2035 486 2093 498
rect 2293 974 2351 986
rect 2293 498 2305 974
rect 2339 498 2351 974
rect 2293 486 2351 498
rect 2551 974 2609 986
rect 2551 498 2563 974
rect 2597 498 2609 974
rect 2551 486 2609 498
rect -2609 238 -2551 250
rect -2609 -238 -2597 238
rect -2563 -238 -2551 238
rect -2609 -250 -2551 -238
rect -2351 238 -2293 250
rect -2351 -238 -2339 238
rect -2305 -238 -2293 238
rect -2351 -250 -2293 -238
rect -2093 238 -2035 250
rect -2093 -238 -2081 238
rect -2047 -238 -2035 238
rect -2093 -250 -2035 -238
rect -1835 238 -1777 250
rect -1835 -238 -1823 238
rect -1789 -238 -1777 238
rect -1835 -250 -1777 -238
rect -1577 238 -1519 250
rect -1577 -238 -1565 238
rect -1531 -238 -1519 238
rect -1577 -250 -1519 -238
rect -1319 238 -1261 250
rect -1319 -238 -1307 238
rect -1273 -238 -1261 238
rect -1319 -250 -1261 -238
rect -1061 238 -1003 250
rect -1061 -238 -1049 238
rect -1015 -238 -1003 238
rect -1061 -250 -1003 -238
rect -803 238 -745 250
rect -803 -238 -791 238
rect -757 -238 -745 238
rect -803 -250 -745 -238
rect -545 238 -487 250
rect -545 -238 -533 238
rect -499 -238 -487 238
rect -545 -250 -487 -238
rect -287 238 -229 250
rect -287 -238 -275 238
rect -241 -238 -229 238
rect -287 -250 -229 -238
rect -29 238 29 250
rect -29 -238 -17 238
rect 17 -238 29 238
rect -29 -250 29 -238
rect 229 238 287 250
rect 229 -238 241 238
rect 275 -238 287 238
rect 229 -250 287 -238
rect 487 238 545 250
rect 487 -238 499 238
rect 533 -238 545 238
rect 487 -250 545 -238
rect 745 238 803 250
rect 745 -238 757 238
rect 791 -238 803 238
rect 745 -250 803 -238
rect 1003 238 1061 250
rect 1003 -238 1015 238
rect 1049 -238 1061 238
rect 1003 -250 1061 -238
rect 1261 238 1319 250
rect 1261 -238 1273 238
rect 1307 -238 1319 238
rect 1261 -250 1319 -238
rect 1519 238 1577 250
rect 1519 -238 1531 238
rect 1565 -238 1577 238
rect 1519 -250 1577 -238
rect 1777 238 1835 250
rect 1777 -238 1789 238
rect 1823 -238 1835 238
rect 1777 -250 1835 -238
rect 2035 238 2093 250
rect 2035 -238 2047 238
rect 2081 -238 2093 238
rect 2035 -250 2093 -238
rect 2293 238 2351 250
rect 2293 -238 2305 238
rect 2339 -238 2351 238
rect 2293 -250 2351 -238
rect 2551 238 2609 250
rect 2551 -238 2563 238
rect 2597 -238 2609 238
rect 2551 -250 2609 -238
rect -2609 -498 -2551 -486
rect -2609 -974 -2597 -498
rect -2563 -974 -2551 -498
rect -2609 -986 -2551 -974
rect -2351 -498 -2293 -486
rect -2351 -974 -2339 -498
rect -2305 -974 -2293 -498
rect -2351 -986 -2293 -974
rect -2093 -498 -2035 -486
rect -2093 -974 -2081 -498
rect -2047 -974 -2035 -498
rect -2093 -986 -2035 -974
rect -1835 -498 -1777 -486
rect -1835 -974 -1823 -498
rect -1789 -974 -1777 -498
rect -1835 -986 -1777 -974
rect -1577 -498 -1519 -486
rect -1577 -974 -1565 -498
rect -1531 -974 -1519 -498
rect -1577 -986 -1519 -974
rect -1319 -498 -1261 -486
rect -1319 -974 -1307 -498
rect -1273 -974 -1261 -498
rect -1319 -986 -1261 -974
rect -1061 -498 -1003 -486
rect -1061 -974 -1049 -498
rect -1015 -974 -1003 -498
rect -1061 -986 -1003 -974
rect -803 -498 -745 -486
rect -803 -974 -791 -498
rect -757 -974 -745 -498
rect -803 -986 -745 -974
rect -545 -498 -487 -486
rect -545 -974 -533 -498
rect -499 -974 -487 -498
rect -545 -986 -487 -974
rect -287 -498 -229 -486
rect -287 -974 -275 -498
rect -241 -974 -229 -498
rect -287 -986 -229 -974
rect -29 -498 29 -486
rect -29 -974 -17 -498
rect 17 -974 29 -498
rect -29 -986 29 -974
rect 229 -498 287 -486
rect 229 -974 241 -498
rect 275 -974 287 -498
rect 229 -986 287 -974
rect 487 -498 545 -486
rect 487 -974 499 -498
rect 533 -974 545 -498
rect 487 -986 545 -974
rect 745 -498 803 -486
rect 745 -974 757 -498
rect 791 -974 803 -498
rect 745 -986 803 -974
rect 1003 -498 1061 -486
rect 1003 -974 1015 -498
rect 1049 -974 1061 -498
rect 1003 -986 1061 -974
rect 1261 -498 1319 -486
rect 1261 -974 1273 -498
rect 1307 -974 1319 -498
rect 1261 -986 1319 -974
rect 1519 -498 1577 -486
rect 1519 -974 1531 -498
rect 1565 -974 1577 -498
rect 1519 -986 1577 -974
rect 1777 -498 1835 -486
rect 1777 -974 1789 -498
rect 1823 -974 1835 -498
rect 1777 -986 1835 -974
rect 2035 -498 2093 -486
rect 2035 -974 2047 -498
rect 2081 -974 2093 -498
rect 2035 -986 2093 -974
rect 2293 -498 2351 -486
rect 2293 -974 2305 -498
rect 2339 -974 2351 -498
rect 2293 -986 2351 -974
rect 2551 -498 2609 -486
rect 2551 -974 2563 -498
rect 2597 -974 2609 -498
rect 2551 -986 2609 -974
rect -2609 -1234 -2551 -1222
rect -2609 -1710 -2597 -1234
rect -2563 -1710 -2551 -1234
rect -2609 -1722 -2551 -1710
rect -2351 -1234 -2293 -1222
rect -2351 -1710 -2339 -1234
rect -2305 -1710 -2293 -1234
rect -2351 -1722 -2293 -1710
rect -2093 -1234 -2035 -1222
rect -2093 -1710 -2081 -1234
rect -2047 -1710 -2035 -1234
rect -2093 -1722 -2035 -1710
rect -1835 -1234 -1777 -1222
rect -1835 -1710 -1823 -1234
rect -1789 -1710 -1777 -1234
rect -1835 -1722 -1777 -1710
rect -1577 -1234 -1519 -1222
rect -1577 -1710 -1565 -1234
rect -1531 -1710 -1519 -1234
rect -1577 -1722 -1519 -1710
rect -1319 -1234 -1261 -1222
rect -1319 -1710 -1307 -1234
rect -1273 -1710 -1261 -1234
rect -1319 -1722 -1261 -1710
rect -1061 -1234 -1003 -1222
rect -1061 -1710 -1049 -1234
rect -1015 -1710 -1003 -1234
rect -1061 -1722 -1003 -1710
rect -803 -1234 -745 -1222
rect -803 -1710 -791 -1234
rect -757 -1710 -745 -1234
rect -803 -1722 -745 -1710
rect -545 -1234 -487 -1222
rect -545 -1710 -533 -1234
rect -499 -1710 -487 -1234
rect -545 -1722 -487 -1710
rect -287 -1234 -229 -1222
rect -287 -1710 -275 -1234
rect -241 -1710 -229 -1234
rect -287 -1722 -229 -1710
rect -29 -1234 29 -1222
rect -29 -1710 -17 -1234
rect 17 -1710 29 -1234
rect -29 -1722 29 -1710
rect 229 -1234 287 -1222
rect 229 -1710 241 -1234
rect 275 -1710 287 -1234
rect 229 -1722 287 -1710
rect 487 -1234 545 -1222
rect 487 -1710 499 -1234
rect 533 -1710 545 -1234
rect 487 -1722 545 -1710
rect 745 -1234 803 -1222
rect 745 -1710 757 -1234
rect 791 -1710 803 -1234
rect 745 -1722 803 -1710
rect 1003 -1234 1061 -1222
rect 1003 -1710 1015 -1234
rect 1049 -1710 1061 -1234
rect 1003 -1722 1061 -1710
rect 1261 -1234 1319 -1222
rect 1261 -1710 1273 -1234
rect 1307 -1710 1319 -1234
rect 1261 -1722 1319 -1710
rect 1519 -1234 1577 -1222
rect 1519 -1710 1531 -1234
rect 1565 -1710 1577 -1234
rect 1519 -1722 1577 -1710
rect 1777 -1234 1835 -1222
rect 1777 -1710 1789 -1234
rect 1823 -1710 1835 -1234
rect 1777 -1722 1835 -1710
rect 2035 -1234 2093 -1222
rect 2035 -1710 2047 -1234
rect 2081 -1710 2093 -1234
rect 2035 -1722 2093 -1710
rect 2293 -1234 2351 -1222
rect 2293 -1710 2305 -1234
rect 2339 -1710 2351 -1234
rect 2293 -1722 2351 -1710
rect 2551 -1234 2609 -1222
rect 2551 -1710 2563 -1234
rect 2597 -1710 2609 -1234
rect 2551 -1722 2609 -1710
rect -2609 -1970 -2551 -1958
rect -2609 -2446 -2597 -1970
rect -2563 -2446 -2551 -1970
rect -2609 -2458 -2551 -2446
rect -2351 -1970 -2293 -1958
rect -2351 -2446 -2339 -1970
rect -2305 -2446 -2293 -1970
rect -2351 -2458 -2293 -2446
rect -2093 -1970 -2035 -1958
rect -2093 -2446 -2081 -1970
rect -2047 -2446 -2035 -1970
rect -2093 -2458 -2035 -2446
rect -1835 -1970 -1777 -1958
rect -1835 -2446 -1823 -1970
rect -1789 -2446 -1777 -1970
rect -1835 -2458 -1777 -2446
rect -1577 -1970 -1519 -1958
rect -1577 -2446 -1565 -1970
rect -1531 -2446 -1519 -1970
rect -1577 -2458 -1519 -2446
rect -1319 -1970 -1261 -1958
rect -1319 -2446 -1307 -1970
rect -1273 -2446 -1261 -1970
rect -1319 -2458 -1261 -2446
rect -1061 -1970 -1003 -1958
rect -1061 -2446 -1049 -1970
rect -1015 -2446 -1003 -1970
rect -1061 -2458 -1003 -2446
rect -803 -1970 -745 -1958
rect -803 -2446 -791 -1970
rect -757 -2446 -745 -1970
rect -803 -2458 -745 -2446
rect -545 -1970 -487 -1958
rect -545 -2446 -533 -1970
rect -499 -2446 -487 -1970
rect -545 -2458 -487 -2446
rect -287 -1970 -229 -1958
rect -287 -2446 -275 -1970
rect -241 -2446 -229 -1970
rect -287 -2458 -229 -2446
rect -29 -1970 29 -1958
rect -29 -2446 -17 -1970
rect 17 -2446 29 -1970
rect -29 -2458 29 -2446
rect 229 -1970 287 -1958
rect 229 -2446 241 -1970
rect 275 -2446 287 -1970
rect 229 -2458 287 -2446
rect 487 -1970 545 -1958
rect 487 -2446 499 -1970
rect 533 -2446 545 -1970
rect 487 -2458 545 -2446
rect 745 -1970 803 -1958
rect 745 -2446 757 -1970
rect 791 -2446 803 -1970
rect 745 -2458 803 -2446
rect 1003 -1970 1061 -1958
rect 1003 -2446 1015 -1970
rect 1049 -2446 1061 -1970
rect 1003 -2458 1061 -2446
rect 1261 -1970 1319 -1958
rect 1261 -2446 1273 -1970
rect 1307 -2446 1319 -1970
rect 1261 -2458 1319 -2446
rect 1519 -1970 1577 -1958
rect 1519 -2446 1531 -1970
rect 1565 -2446 1577 -1970
rect 1519 -2458 1577 -2446
rect 1777 -1970 1835 -1958
rect 1777 -2446 1789 -1970
rect 1823 -2446 1835 -1970
rect 1777 -2458 1835 -2446
rect 2035 -1970 2093 -1958
rect 2035 -2446 2047 -1970
rect 2081 -2446 2093 -1970
rect 2035 -2458 2093 -2446
rect 2293 -1970 2351 -1958
rect 2293 -2446 2305 -1970
rect 2339 -2446 2351 -1970
rect 2293 -2458 2351 -2446
rect 2551 -1970 2609 -1958
rect 2551 -2446 2563 -1970
rect 2597 -2446 2609 -1970
rect 2551 -2458 2609 -2446
<< pdiffc >>
rect -2597 1970 -2563 2446
rect -2339 1970 -2305 2446
rect -2081 1970 -2047 2446
rect -1823 1970 -1789 2446
rect -1565 1970 -1531 2446
rect -1307 1970 -1273 2446
rect -1049 1970 -1015 2446
rect -791 1970 -757 2446
rect -533 1970 -499 2446
rect -275 1970 -241 2446
rect -17 1970 17 2446
rect 241 1970 275 2446
rect 499 1970 533 2446
rect 757 1970 791 2446
rect 1015 1970 1049 2446
rect 1273 1970 1307 2446
rect 1531 1970 1565 2446
rect 1789 1970 1823 2446
rect 2047 1970 2081 2446
rect 2305 1970 2339 2446
rect 2563 1970 2597 2446
rect -2597 1234 -2563 1710
rect -2339 1234 -2305 1710
rect -2081 1234 -2047 1710
rect -1823 1234 -1789 1710
rect -1565 1234 -1531 1710
rect -1307 1234 -1273 1710
rect -1049 1234 -1015 1710
rect -791 1234 -757 1710
rect -533 1234 -499 1710
rect -275 1234 -241 1710
rect -17 1234 17 1710
rect 241 1234 275 1710
rect 499 1234 533 1710
rect 757 1234 791 1710
rect 1015 1234 1049 1710
rect 1273 1234 1307 1710
rect 1531 1234 1565 1710
rect 1789 1234 1823 1710
rect 2047 1234 2081 1710
rect 2305 1234 2339 1710
rect 2563 1234 2597 1710
rect -2597 498 -2563 974
rect -2339 498 -2305 974
rect -2081 498 -2047 974
rect -1823 498 -1789 974
rect -1565 498 -1531 974
rect -1307 498 -1273 974
rect -1049 498 -1015 974
rect -791 498 -757 974
rect -533 498 -499 974
rect -275 498 -241 974
rect -17 498 17 974
rect 241 498 275 974
rect 499 498 533 974
rect 757 498 791 974
rect 1015 498 1049 974
rect 1273 498 1307 974
rect 1531 498 1565 974
rect 1789 498 1823 974
rect 2047 498 2081 974
rect 2305 498 2339 974
rect 2563 498 2597 974
rect -2597 -238 -2563 238
rect -2339 -238 -2305 238
rect -2081 -238 -2047 238
rect -1823 -238 -1789 238
rect -1565 -238 -1531 238
rect -1307 -238 -1273 238
rect -1049 -238 -1015 238
rect -791 -238 -757 238
rect -533 -238 -499 238
rect -275 -238 -241 238
rect -17 -238 17 238
rect 241 -238 275 238
rect 499 -238 533 238
rect 757 -238 791 238
rect 1015 -238 1049 238
rect 1273 -238 1307 238
rect 1531 -238 1565 238
rect 1789 -238 1823 238
rect 2047 -238 2081 238
rect 2305 -238 2339 238
rect 2563 -238 2597 238
rect -2597 -974 -2563 -498
rect -2339 -974 -2305 -498
rect -2081 -974 -2047 -498
rect -1823 -974 -1789 -498
rect -1565 -974 -1531 -498
rect -1307 -974 -1273 -498
rect -1049 -974 -1015 -498
rect -791 -974 -757 -498
rect -533 -974 -499 -498
rect -275 -974 -241 -498
rect -17 -974 17 -498
rect 241 -974 275 -498
rect 499 -974 533 -498
rect 757 -974 791 -498
rect 1015 -974 1049 -498
rect 1273 -974 1307 -498
rect 1531 -974 1565 -498
rect 1789 -974 1823 -498
rect 2047 -974 2081 -498
rect 2305 -974 2339 -498
rect 2563 -974 2597 -498
rect -2597 -1710 -2563 -1234
rect -2339 -1710 -2305 -1234
rect -2081 -1710 -2047 -1234
rect -1823 -1710 -1789 -1234
rect -1565 -1710 -1531 -1234
rect -1307 -1710 -1273 -1234
rect -1049 -1710 -1015 -1234
rect -791 -1710 -757 -1234
rect -533 -1710 -499 -1234
rect -275 -1710 -241 -1234
rect -17 -1710 17 -1234
rect 241 -1710 275 -1234
rect 499 -1710 533 -1234
rect 757 -1710 791 -1234
rect 1015 -1710 1049 -1234
rect 1273 -1710 1307 -1234
rect 1531 -1710 1565 -1234
rect 1789 -1710 1823 -1234
rect 2047 -1710 2081 -1234
rect 2305 -1710 2339 -1234
rect 2563 -1710 2597 -1234
rect -2597 -2446 -2563 -1970
rect -2339 -2446 -2305 -1970
rect -2081 -2446 -2047 -1970
rect -1823 -2446 -1789 -1970
rect -1565 -2446 -1531 -1970
rect -1307 -2446 -1273 -1970
rect -1049 -2446 -1015 -1970
rect -791 -2446 -757 -1970
rect -533 -2446 -499 -1970
rect -275 -2446 -241 -1970
rect -17 -2446 17 -1970
rect 241 -2446 275 -1970
rect 499 -2446 533 -1970
rect 757 -2446 791 -1970
rect 1015 -2446 1049 -1970
rect 1273 -2446 1307 -1970
rect 1531 -2446 1565 -1970
rect 1789 -2446 1823 -1970
rect 2047 -2446 2081 -1970
rect 2305 -2446 2339 -1970
rect 2563 -2446 2597 -1970
<< nsubdiff >>
rect -2711 2607 -2615 2641
rect 2615 2607 2711 2641
rect -2711 2545 -2677 2607
rect 2677 2545 2711 2607
rect -2711 -2607 -2677 -2545
rect 2677 -2607 2711 -2545
rect -2711 -2641 -2615 -2607
rect 2615 -2641 2711 -2607
<< nsubdiffcont >>
rect -2615 2607 2615 2641
rect -2711 -2545 -2677 2545
rect 2677 -2545 2711 2545
rect -2615 -2641 2615 -2607
<< poly >>
rect -2551 2539 -2351 2555
rect -2551 2505 -2535 2539
rect -2367 2505 -2351 2539
rect -2551 2458 -2351 2505
rect -2293 2539 -2093 2555
rect -2293 2505 -2277 2539
rect -2109 2505 -2093 2539
rect -2293 2458 -2093 2505
rect -2035 2539 -1835 2555
rect -2035 2505 -2019 2539
rect -1851 2505 -1835 2539
rect -2035 2458 -1835 2505
rect -1777 2539 -1577 2555
rect -1777 2505 -1761 2539
rect -1593 2505 -1577 2539
rect -1777 2458 -1577 2505
rect -1519 2539 -1319 2555
rect -1519 2505 -1503 2539
rect -1335 2505 -1319 2539
rect -1519 2458 -1319 2505
rect -1261 2539 -1061 2555
rect -1261 2505 -1245 2539
rect -1077 2505 -1061 2539
rect -1261 2458 -1061 2505
rect -1003 2539 -803 2555
rect -1003 2505 -987 2539
rect -819 2505 -803 2539
rect -1003 2458 -803 2505
rect -745 2539 -545 2555
rect -745 2505 -729 2539
rect -561 2505 -545 2539
rect -745 2458 -545 2505
rect -487 2539 -287 2555
rect -487 2505 -471 2539
rect -303 2505 -287 2539
rect -487 2458 -287 2505
rect -229 2539 -29 2555
rect -229 2505 -213 2539
rect -45 2505 -29 2539
rect -229 2458 -29 2505
rect 29 2539 229 2555
rect 29 2505 45 2539
rect 213 2505 229 2539
rect 29 2458 229 2505
rect 287 2539 487 2555
rect 287 2505 303 2539
rect 471 2505 487 2539
rect 287 2458 487 2505
rect 545 2539 745 2555
rect 545 2505 561 2539
rect 729 2505 745 2539
rect 545 2458 745 2505
rect 803 2539 1003 2555
rect 803 2505 819 2539
rect 987 2505 1003 2539
rect 803 2458 1003 2505
rect 1061 2539 1261 2555
rect 1061 2505 1077 2539
rect 1245 2505 1261 2539
rect 1061 2458 1261 2505
rect 1319 2539 1519 2555
rect 1319 2505 1335 2539
rect 1503 2505 1519 2539
rect 1319 2458 1519 2505
rect 1577 2539 1777 2555
rect 1577 2505 1593 2539
rect 1761 2505 1777 2539
rect 1577 2458 1777 2505
rect 1835 2539 2035 2555
rect 1835 2505 1851 2539
rect 2019 2505 2035 2539
rect 1835 2458 2035 2505
rect 2093 2539 2293 2555
rect 2093 2505 2109 2539
rect 2277 2505 2293 2539
rect 2093 2458 2293 2505
rect 2351 2539 2551 2555
rect 2351 2505 2367 2539
rect 2535 2505 2551 2539
rect 2351 2458 2551 2505
rect -2551 1911 -2351 1958
rect -2551 1877 -2535 1911
rect -2367 1877 -2351 1911
rect -2551 1861 -2351 1877
rect -2293 1911 -2093 1958
rect -2293 1877 -2277 1911
rect -2109 1877 -2093 1911
rect -2293 1861 -2093 1877
rect -2035 1911 -1835 1958
rect -2035 1877 -2019 1911
rect -1851 1877 -1835 1911
rect -2035 1861 -1835 1877
rect -1777 1911 -1577 1958
rect -1777 1877 -1761 1911
rect -1593 1877 -1577 1911
rect -1777 1861 -1577 1877
rect -1519 1911 -1319 1958
rect -1519 1877 -1503 1911
rect -1335 1877 -1319 1911
rect -1519 1861 -1319 1877
rect -1261 1911 -1061 1958
rect -1261 1877 -1245 1911
rect -1077 1877 -1061 1911
rect -1261 1861 -1061 1877
rect -1003 1911 -803 1958
rect -1003 1877 -987 1911
rect -819 1877 -803 1911
rect -1003 1861 -803 1877
rect -745 1911 -545 1958
rect -745 1877 -729 1911
rect -561 1877 -545 1911
rect -745 1861 -545 1877
rect -487 1911 -287 1958
rect -487 1877 -471 1911
rect -303 1877 -287 1911
rect -487 1861 -287 1877
rect -229 1911 -29 1958
rect -229 1877 -213 1911
rect -45 1877 -29 1911
rect -229 1861 -29 1877
rect 29 1911 229 1958
rect 29 1877 45 1911
rect 213 1877 229 1911
rect 29 1861 229 1877
rect 287 1911 487 1958
rect 287 1877 303 1911
rect 471 1877 487 1911
rect 287 1861 487 1877
rect 545 1911 745 1958
rect 545 1877 561 1911
rect 729 1877 745 1911
rect 545 1861 745 1877
rect 803 1911 1003 1958
rect 803 1877 819 1911
rect 987 1877 1003 1911
rect 803 1861 1003 1877
rect 1061 1911 1261 1958
rect 1061 1877 1077 1911
rect 1245 1877 1261 1911
rect 1061 1861 1261 1877
rect 1319 1911 1519 1958
rect 1319 1877 1335 1911
rect 1503 1877 1519 1911
rect 1319 1861 1519 1877
rect 1577 1911 1777 1958
rect 1577 1877 1593 1911
rect 1761 1877 1777 1911
rect 1577 1861 1777 1877
rect 1835 1911 2035 1958
rect 1835 1877 1851 1911
rect 2019 1877 2035 1911
rect 1835 1861 2035 1877
rect 2093 1911 2293 1958
rect 2093 1877 2109 1911
rect 2277 1877 2293 1911
rect 2093 1861 2293 1877
rect 2351 1911 2551 1958
rect 2351 1877 2367 1911
rect 2535 1877 2551 1911
rect 2351 1861 2551 1877
rect -2551 1803 -2351 1819
rect -2551 1769 -2535 1803
rect -2367 1769 -2351 1803
rect -2551 1722 -2351 1769
rect -2293 1803 -2093 1819
rect -2293 1769 -2277 1803
rect -2109 1769 -2093 1803
rect -2293 1722 -2093 1769
rect -2035 1803 -1835 1819
rect -2035 1769 -2019 1803
rect -1851 1769 -1835 1803
rect -2035 1722 -1835 1769
rect -1777 1803 -1577 1819
rect -1777 1769 -1761 1803
rect -1593 1769 -1577 1803
rect -1777 1722 -1577 1769
rect -1519 1803 -1319 1819
rect -1519 1769 -1503 1803
rect -1335 1769 -1319 1803
rect -1519 1722 -1319 1769
rect -1261 1803 -1061 1819
rect -1261 1769 -1245 1803
rect -1077 1769 -1061 1803
rect -1261 1722 -1061 1769
rect -1003 1803 -803 1819
rect -1003 1769 -987 1803
rect -819 1769 -803 1803
rect -1003 1722 -803 1769
rect -745 1803 -545 1819
rect -745 1769 -729 1803
rect -561 1769 -545 1803
rect -745 1722 -545 1769
rect -487 1803 -287 1819
rect -487 1769 -471 1803
rect -303 1769 -287 1803
rect -487 1722 -287 1769
rect -229 1803 -29 1819
rect -229 1769 -213 1803
rect -45 1769 -29 1803
rect -229 1722 -29 1769
rect 29 1803 229 1819
rect 29 1769 45 1803
rect 213 1769 229 1803
rect 29 1722 229 1769
rect 287 1803 487 1819
rect 287 1769 303 1803
rect 471 1769 487 1803
rect 287 1722 487 1769
rect 545 1803 745 1819
rect 545 1769 561 1803
rect 729 1769 745 1803
rect 545 1722 745 1769
rect 803 1803 1003 1819
rect 803 1769 819 1803
rect 987 1769 1003 1803
rect 803 1722 1003 1769
rect 1061 1803 1261 1819
rect 1061 1769 1077 1803
rect 1245 1769 1261 1803
rect 1061 1722 1261 1769
rect 1319 1803 1519 1819
rect 1319 1769 1335 1803
rect 1503 1769 1519 1803
rect 1319 1722 1519 1769
rect 1577 1803 1777 1819
rect 1577 1769 1593 1803
rect 1761 1769 1777 1803
rect 1577 1722 1777 1769
rect 1835 1803 2035 1819
rect 1835 1769 1851 1803
rect 2019 1769 2035 1803
rect 1835 1722 2035 1769
rect 2093 1803 2293 1819
rect 2093 1769 2109 1803
rect 2277 1769 2293 1803
rect 2093 1722 2293 1769
rect 2351 1803 2551 1819
rect 2351 1769 2367 1803
rect 2535 1769 2551 1803
rect 2351 1722 2551 1769
rect -2551 1175 -2351 1222
rect -2551 1141 -2535 1175
rect -2367 1141 -2351 1175
rect -2551 1125 -2351 1141
rect -2293 1175 -2093 1222
rect -2293 1141 -2277 1175
rect -2109 1141 -2093 1175
rect -2293 1125 -2093 1141
rect -2035 1175 -1835 1222
rect -2035 1141 -2019 1175
rect -1851 1141 -1835 1175
rect -2035 1125 -1835 1141
rect -1777 1175 -1577 1222
rect -1777 1141 -1761 1175
rect -1593 1141 -1577 1175
rect -1777 1125 -1577 1141
rect -1519 1175 -1319 1222
rect -1519 1141 -1503 1175
rect -1335 1141 -1319 1175
rect -1519 1125 -1319 1141
rect -1261 1175 -1061 1222
rect -1261 1141 -1245 1175
rect -1077 1141 -1061 1175
rect -1261 1125 -1061 1141
rect -1003 1175 -803 1222
rect -1003 1141 -987 1175
rect -819 1141 -803 1175
rect -1003 1125 -803 1141
rect -745 1175 -545 1222
rect -745 1141 -729 1175
rect -561 1141 -545 1175
rect -745 1125 -545 1141
rect -487 1175 -287 1222
rect -487 1141 -471 1175
rect -303 1141 -287 1175
rect -487 1125 -287 1141
rect -229 1175 -29 1222
rect -229 1141 -213 1175
rect -45 1141 -29 1175
rect -229 1125 -29 1141
rect 29 1175 229 1222
rect 29 1141 45 1175
rect 213 1141 229 1175
rect 29 1125 229 1141
rect 287 1175 487 1222
rect 287 1141 303 1175
rect 471 1141 487 1175
rect 287 1125 487 1141
rect 545 1175 745 1222
rect 545 1141 561 1175
rect 729 1141 745 1175
rect 545 1125 745 1141
rect 803 1175 1003 1222
rect 803 1141 819 1175
rect 987 1141 1003 1175
rect 803 1125 1003 1141
rect 1061 1175 1261 1222
rect 1061 1141 1077 1175
rect 1245 1141 1261 1175
rect 1061 1125 1261 1141
rect 1319 1175 1519 1222
rect 1319 1141 1335 1175
rect 1503 1141 1519 1175
rect 1319 1125 1519 1141
rect 1577 1175 1777 1222
rect 1577 1141 1593 1175
rect 1761 1141 1777 1175
rect 1577 1125 1777 1141
rect 1835 1175 2035 1222
rect 1835 1141 1851 1175
rect 2019 1141 2035 1175
rect 1835 1125 2035 1141
rect 2093 1175 2293 1222
rect 2093 1141 2109 1175
rect 2277 1141 2293 1175
rect 2093 1125 2293 1141
rect 2351 1175 2551 1222
rect 2351 1141 2367 1175
rect 2535 1141 2551 1175
rect 2351 1125 2551 1141
rect -2551 1067 -2351 1083
rect -2551 1033 -2535 1067
rect -2367 1033 -2351 1067
rect -2551 986 -2351 1033
rect -2293 1067 -2093 1083
rect -2293 1033 -2277 1067
rect -2109 1033 -2093 1067
rect -2293 986 -2093 1033
rect -2035 1067 -1835 1083
rect -2035 1033 -2019 1067
rect -1851 1033 -1835 1067
rect -2035 986 -1835 1033
rect -1777 1067 -1577 1083
rect -1777 1033 -1761 1067
rect -1593 1033 -1577 1067
rect -1777 986 -1577 1033
rect -1519 1067 -1319 1083
rect -1519 1033 -1503 1067
rect -1335 1033 -1319 1067
rect -1519 986 -1319 1033
rect -1261 1067 -1061 1083
rect -1261 1033 -1245 1067
rect -1077 1033 -1061 1067
rect -1261 986 -1061 1033
rect -1003 1067 -803 1083
rect -1003 1033 -987 1067
rect -819 1033 -803 1067
rect -1003 986 -803 1033
rect -745 1067 -545 1083
rect -745 1033 -729 1067
rect -561 1033 -545 1067
rect -745 986 -545 1033
rect -487 1067 -287 1083
rect -487 1033 -471 1067
rect -303 1033 -287 1067
rect -487 986 -287 1033
rect -229 1067 -29 1083
rect -229 1033 -213 1067
rect -45 1033 -29 1067
rect -229 986 -29 1033
rect 29 1067 229 1083
rect 29 1033 45 1067
rect 213 1033 229 1067
rect 29 986 229 1033
rect 287 1067 487 1083
rect 287 1033 303 1067
rect 471 1033 487 1067
rect 287 986 487 1033
rect 545 1067 745 1083
rect 545 1033 561 1067
rect 729 1033 745 1067
rect 545 986 745 1033
rect 803 1067 1003 1083
rect 803 1033 819 1067
rect 987 1033 1003 1067
rect 803 986 1003 1033
rect 1061 1067 1261 1083
rect 1061 1033 1077 1067
rect 1245 1033 1261 1067
rect 1061 986 1261 1033
rect 1319 1067 1519 1083
rect 1319 1033 1335 1067
rect 1503 1033 1519 1067
rect 1319 986 1519 1033
rect 1577 1067 1777 1083
rect 1577 1033 1593 1067
rect 1761 1033 1777 1067
rect 1577 986 1777 1033
rect 1835 1067 2035 1083
rect 1835 1033 1851 1067
rect 2019 1033 2035 1067
rect 1835 986 2035 1033
rect 2093 1067 2293 1083
rect 2093 1033 2109 1067
rect 2277 1033 2293 1067
rect 2093 986 2293 1033
rect 2351 1067 2551 1083
rect 2351 1033 2367 1067
rect 2535 1033 2551 1067
rect 2351 986 2551 1033
rect -2551 439 -2351 486
rect -2551 405 -2535 439
rect -2367 405 -2351 439
rect -2551 389 -2351 405
rect -2293 439 -2093 486
rect -2293 405 -2277 439
rect -2109 405 -2093 439
rect -2293 389 -2093 405
rect -2035 439 -1835 486
rect -2035 405 -2019 439
rect -1851 405 -1835 439
rect -2035 389 -1835 405
rect -1777 439 -1577 486
rect -1777 405 -1761 439
rect -1593 405 -1577 439
rect -1777 389 -1577 405
rect -1519 439 -1319 486
rect -1519 405 -1503 439
rect -1335 405 -1319 439
rect -1519 389 -1319 405
rect -1261 439 -1061 486
rect -1261 405 -1245 439
rect -1077 405 -1061 439
rect -1261 389 -1061 405
rect -1003 439 -803 486
rect -1003 405 -987 439
rect -819 405 -803 439
rect -1003 389 -803 405
rect -745 439 -545 486
rect -745 405 -729 439
rect -561 405 -545 439
rect -745 389 -545 405
rect -487 439 -287 486
rect -487 405 -471 439
rect -303 405 -287 439
rect -487 389 -287 405
rect -229 439 -29 486
rect -229 405 -213 439
rect -45 405 -29 439
rect -229 389 -29 405
rect 29 439 229 486
rect 29 405 45 439
rect 213 405 229 439
rect 29 389 229 405
rect 287 439 487 486
rect 287 405 303 439
rect 471 405 487 439
rect 287 389 487 405
rect 545 439 745 486
rect 545 405 561 439
rect 729 405 745 439
rect 545 389 745 405
rect 803 439 1003 486
rect 803 405 819 439
rect 987 405 1003 439
rect 803 389 1003 405
rect 1061 439 1261 486
rect 1061 405 1077 439
rect 1245 405 1261 439
rect 1061 389 1261 405
rect 1319 439 1519 486
rect 1319 405 1335 439
rect 1503 405 1519 439
rect 1319 389 1519 405
rect 1577 439 1777 486
rect 1577 405 1593 439
rect 1761 405 1777 439
rect 1577 389 1777 405
rect 1835 439 2035 486
rect 1835 405 1851 439
rect 2019 405 2035 439
rect 1835 389 2035 405
rect 2093 439 2293 486
rect 2093 405 2109 439
rect 2277 405 2293 439
rect 2093 389 2293 405
rect 2351 439 2551 486
rect 2351 405 2367 439
rect 2535 405 2551 439
rect 2351 389 2551 405
rect -2551 331 -2351 347
rect -2551 297 -2535 331
rect -2367 297 -2351 331
rect -2551 250 -2351 297
rect -2293 331 -2093 347
rect -2293 297 -2277 331
rect -2109 297 -2093 331
rect -2293 250 -2093 297
rect -2035 331 -1835 347
rect -2035 297 -2019 331
rect -1851 297 -1835 331
rect -2035 250 -1835 297
rect -1777 331 -1577 347
rect -1777 297 -1761 331
rect -1593 297 -1577 331
rect -1777 250 -1577 297
rect -1519 331 -1319 347
rect -1519 297 -1503 331
rect -1335 297 -1319 331
rect -1519 250 -1319 297
rect -1261 331 -1061 347
rect -1261 297 -1245 331
rect -1077 297 -1061 331
rect -1261 250 -1061 297
rect -1003 331 -803 347
rect -1003 297 -987 331
rect -819 297 -803 331
rect -1003 250 -803 297
rect -745 331 -545 347
rect -745 297 -729 331
rect -561 297 -545 331
rect -745 250 -545 297
rect -487 331 -287 347
rect -487 297 -471 331
rect -303 297 -287 331
rect -487 250 -287 297
rect -229 331 -29 347
rect -229 297 -213 331
rect -45 297 -29 331
rect -229 250 -29 297
rect 29 331 229 347
rect 29 297 45 331
rect 213 297 229 331
rect 29 250 229 297
rect 287 331 487 347
rect 287 297 303 331
rect 471 297 487 331
rect 287 250 487 297
rect 545 331 745 347
rect 545 297 561 331
rect 729 297 745 331
rect 545 250 745 297
rect 803 331 1003 347
rect 803 297 819 331
rect 987 297 1003 331
rect 803 250 1003 297
rect 1061 331 1261 347
rect 1061 297 1077 331
rect 1245 297 1261 331
rect 1061 250 1261 297
rect 1319 331 1519 347
rect 1319 297 1335 331
rect 1503 297 1519 331
rect 1319 250 1519 297
rect 1577 331 1777 347
rect 1577 297 1593 331
rect 1761 297 1777 331
rect 1577 250 1777 297
rect 1835 331 2035 347
rect 1835 297 1851 331
rect 2019 297 2035 331
rect 1835 250 2035 297
rect 2093 331 2293 347
rect 2093 297 2109 331
rect 2277 297 2293 331
rect 2093 250 2293 297
rect 2351 331 2551 347
rect 2351 297 2367 331
rect 2535 297 2551 331
rect 2351 250 2551 297
rect -2551 -297 -2351 -250
rect -2551 -331 -2535 -297
rect -2367 -331 -2351 -297
rect -2551 -347 -2351 -331
rect -2293 -297 -2093 -250
rect -2293 -331 -2277 -297
rect -2109 -331 -2093 -297
rect -2293 -347 -2093 -331
rect -2035 -297 -1835 -250
rect -2035 -331 -2019 -297
rect -1851 -331 -1835 -297
rect -2035 -347 -1835 -331
rect -1777 -297 -1577 -250
rect -1777 -331 -1761 -297
rect -1593 -331 -1577 -297
rect -1777 -347 -1577 -331
rect -1519 -297 -1319 -250
rect -1519 -331 -1503 -297
rect -1335 -331 -1319 -297
rect -1519 -347 -1319 -331
rect -1261 -297 -1061 -250
rect -1261 -331 -1245 -297
rect -1077 -331 -1061 -297
rect -1261 -347 -1061 -331
rect -1003 -297 -803 -250
rect -1003 -331 -987 -297
rect -819 -331 -803 -297
rect -1003 -347 -803 -331
rect -745 -297 -545 -250
rect -745 -331 -729 -297
rect -561 -331 -545 -297
rect -745 -347 -545 -331
rect -487 -297 -287 -250
rect -487 -331 -471 -297
rect -303 -331 -287 -297
rect -487 -347 -287 -331
rect -229 -297 -29 -250
rect -229 -331 -213 -297
rect -45 -331 -29 -297
rect -229 -347 -29 -331
rect 29 -297 229 -250
rect 29 -331 45 -297
rect 213 -331 229 -297
rect 29 -347 229 -331
rect 287 -297 487 -250
rect 287 -331 303 -297
rect 471 -331 487 -297
rect 287 -347 487 -331
rect 545 -297 745 -250
rect 545 -331 561 -297
rect 729 -331 745 -297
rect 545 -347 745 -331
rect 803 -297 1003 -250
rect 803 -331 819 -297
rect 987 -331 1003 -297
rect 803 -347 1003 -331
rect 1061 -297 1261 -250
rect 1061 -331 1077 -297
rect 1245 -331 1261 -297
rect 1061 -347 1261 -331
rect 1319 -297 1519 -250
rect 1319 -331 1335 -297
rect 1503 -331 1519 -297
rect 1319 -347 1519 -331
rect 1577 -297 1777 -250
rect 1577 -331 1593 -297
rect 1761 -331 1777 -297
rect 1577 -347 1777 -331
rect 1835 -297 2035 -250
rect 1835 -331 1851 -297
rect 2019 -331 2035 -297
rect 1835 -347 2035 -331
rect 2093 -297 2293 -250
rect 2093 -331 2109 -297
rect 2277 -331 2293 -297
rect 2093 -347 2293 -331
rect 2351 -297 2551 -250
rect 2351 -331 2367 -297
rect 2535 -331 2551 -297
rect 2351 -347 2551 -331
rect -2551 -405 -2351 -389
rect -2551 -439 -2535 -405
rect -2367 -439 -2351 -405
rect -2551 -486 -2351 -439
rect -2293 -405 -2093 -389
rect -2293 -439 -2277 -405
rect -2109 -439 -2093 -405
rect -2293 -486 -2093 -439
rect -2035 -405 -1835 -389
rect -2035 -439 -2019 -405
rect -1851 -439 -1835 -405
rect -2035 -486 -1835 -439
rect -1777 -405 -1577 -389
rect -1777 -439 -1761 -405
rect -1593 -439 -1577 -405
rect -1777 -486 -1577 -439
rect -1519 -405 -1319 -389
rect -1519 -439 -1503 -405
rect -1335 -439 -1319 -405
rect -1519 -486 -1319 -439
rect -1261 -405 -1061 -389
rect -1261 -439 -1245 -405
rect -1077 -439 -1061 -405
rect -1261 -486 -1061 -439
rect -1003 -405 -803 -389
rect -1003 -439 -987 -405
rect -819 -439 -803 -405
rect -1003 -486 -803 -439
rect -745 -405 -545 -389
rect -745 -439 -729 -405
rect -561 -439 -545 -405
rect -745 -486 -545 -439
rect -487 -405 -287 -389
rect -487 -439 -471 -405
rect -303 -439 -287 -405
rect -487 -486 -287 -439
rect -229 -405 -29 -389
rect -229 -439 -213 -405
rect -45 -439 -29 -405
rect -229 -486 -29 -439
rect 29 -405 229 -389
rect 29 -439 45 -405
rect 213 -439 229 -405
rect 29 -486 229 -439
rect 287 -405 487 -389
rect 287 -439 303 -405
rect 471 -439 487 -405
rect 287 -486 487 -439
rect 545 -405 745 -389
rect 545 -439 561 -405
rect 729 -439 745 -405
rect 545 -486 745 -439
rect 803 -405 1003 -389
rect 803 -439 819 -405
rect 987 -439 1003 -405
rect 803 -486 1003 -439
rect 1061 -405 1261 -389
rect 1061 -439 1077 -405
rect 1245 -439 1261 -405
rect 1061 -486 1261 -439
rect 1319 -405 1519 -389
rect 1319 -439 1335 -405
rect 1503 -439 1519 -405
rect 1319 -486 1519 -439
rect 1577 -405 1777 -389
rect 1577 -439 1593 -405
rect 1761 -439 1777 -405
rect 1577 -486 1777 -439
rect 1835 -405 2035 -389
rect 1835 -439 1851 -405
rect 2019 -439 2035 -405
rect 1835 -486 2035 -439
rect 2093 -405 2293 -389
rect 2093 -439 2109 -405
rect 2277 -439 2293 -405
rect 2093 -486 2293 -439
rect 2351 -405 2551 -389
rect 2351 -439 2367 -405
rect 2535 -439 2551 -405
rect 2351 -486 2551 -439
rect -2551 -1033 -2351 -986
rect -2551 -1067 -2535 -1033
rect -2367 -1067 -2351 -1033
rect -2551 -1083 -2351 -1067
rect -2293 -1033 -2093 -986
rect -2293 -1067 -2277 -1033
rect -2109 -1067 -2093 -1033
rect -2293 -1083 -2093 -1067
rect -2035 -1033 -1835 -986
rect -2035 -1067 -2019 -1033
rect -1851 -1067 -1835 -1033
rect -2035 -1083 -1835 -1067
rect -1777 -1033 -1577 -986
rect -1777 -1067 -1761 -1033
rect -1593 -1067 -1577 -1033
rect -1777 -1083 -1577 -1067
rect -1519 -1033 -1319 -986
rect -1519 -1067 -1503 -1033
rect -1335 -1067 -1319 -1033
rect -1519 -1083 -1319 -1067
rect -1261 -1033 -1061 -986
rect -1261 -1067 -1245 -1033
rect -1077 -1067 -1061 -1033
rect -1261 -1083 -1061 -1067
rect -1003 -1033 -803 -986
rect -1003 -1067 -987 -1033
rect -819 -1067 -803 -1033
rect -1003 -1083 -803 -1067
rect -745 -1033 -545 -986
rect -745 -1067 -729 -1033
rect -561 -1067 -545 -1033
rect -745 -1083 -545 -1067
rect -487 -1033 -287 -986
rect -487 -1067 -471 -1033
rect -303 -1067 -287 -1033
rect -487 -1083 -287 -1067
rect -229 -1033 -29 -986
rect -229 -1067 -213 -1033
rect -45 -1067 -29 -1033
rect -229 -1083 -29 -1067
rect 29 -1033 229 -986
rect 29 -1067 45 -1033
rect 213 -1067 229 -1033
rect 29 -1083 229 -1067
rect 287 -1033 487 -986
rect 287 -1067 303 -1033
rect 471 -1067 487 -1033
rect 287 -1083 487 -1067
rect 545 -1033 745 -986
rect 545 -1067 561 -1033
rect 729 -1067 745 -1033
rect 545 -1083 745 -1067
rect 803 -1033 1003 -986
rect 803 -1067 819 -1033
rect 987 -1067 1003 -1033
rect 803 -1083 1003 -1067
rect 1061 -1033 1261 -986
rect 1061 -1067 1077 -1033
rect 1245 -1067 1261 -1033
rect 1061 -1083 1261 -1067
rect 1319 -1033 1519 -986
rect 1319 -1067 1335 -1033
rect 1503 -1067 1519 -1033
rect 1319 -1083 1519 -1067
rect 1577 -1033 1777 -986
rect 1577 -1067 1593 -1033
rect 1761 -1067 1777 -1033
rect 1577 -1083 1777 -1067
rect 1835 -1033 2035 -986
rect 1835 -1067 1851 -1033
rect 2019 -1067 2035 -1033
rect 1835 -1083 2035 -1067
rect 2093 -1033 2293 -986
rect 2093 -1067 2109 -1033
rect 2277 -1067 2293 -1033
rect 2093 -1083 2293 -1067
rect 2351 -1033 2551 -986
rect 2351 -1067 2367 -1033
rect 2535 -1067 2551 -1033
rect 2351 -1083 2551 -1067
rect -2551 -1141 -2351 -1125
rect -2551 -1175 -2535 -1141
rect -2367 -1175 -2351 -1141
rect -2551 -1222 -2351 -1175
rect -2293 -1141 -2093 -1125
rect -2293 -1175 -2277 -1141
rect -2109 -1175 -2093 -1141
rect -2293 -1222 -2093 -1175
rect -2035 -1141 -1835 -1125
rect -2035 -1175 -2019 -1141
rect -1851 -1175 -1835 -1141
rect -2035 -1222 -1835 -1175
rect -1777 -1141 -1577 -1125
rect -1777 -1175 -1761 -1141
rect -1593 -1175 -1577 -1141
rect -1777 -1222 -1577 -1175
rect -1519 -1141 -1319 -1125
rect -1519 -1175 -1503 -1141
rect -1335 -1175 -1319 -1141
rect -1519 -1222 -1319 -1175
rect -1261 -1141 -1061 -1125
rect -1261 -1175 -1245 -1141
rect -1077 -1175 -1061 -1141
rect -1261 -1222 -1061 -1175
rect -1003 -1141 -803 -1125
rect -1003 -1175 -987 -1141
rect -819 -1175 -803 -1141
rect -1003 -1222 -803 -1175
rect -745 -1141 -545 -1125
rect -745 -1175 -729 -1141
rect -561 -1175 -545 -1141
rect -745 -1222 -545 -1175
rect -487 -1141 -287 -1125
rect -487 -1175 -471 -1141
rect -303 -1175 -287 -1141
rect -487 -1222 -287 -1175
rect -229 -1141 -29 -1125
rect -229 -1175 -213 -1141
rect -45 -1175 -29 -1141
rect -229 -1222 -29 -1175
rect 29 -1141 229 -1125
rect 29 -1175 45 -1141
rect 213 -1175 229 -1141
rect 29 -1222 229 -1175
rect 287 -1141 487 -1125
rect 287 -1175 303 -1141
rect 471 -1175 487 -1141
rect 287 -1222 487 -1175
rect 545 -1141 745 -1125
rect 545 -1175 561 -1141
rect 729 -1175 745 -1141
rect 545 -1222 745 -1175
rect 803 -1141 1003 -1125
rect 803 -1175 819 -1141
rect 987 -1175 1003 -1141
rect 803 -1222 1003 -1175
rect 1061 -1141 1261 -1125
rect 1061 -1175 1077 -1141
rect 1245 -1175 1261 -1141
rect 1061 -1222 1261 -1175
rect 1319 -1141 1519 -1125
rect 1319 -1175 1335 -1141
rect 1503 -1175 1519 -1141
rect 1319 -1222 1519 -1175
rect 1577 -1141 1777 -1125
rect 1577 -1175 1593 -1141
rect 1761 -1175 1777 -1141
rect 1577 -1222 1777 -1175
rect 1835 -1141 2035 -1125
rect 1835 -1175 1851 -1141
rect 2019 -1175 2035 -1141
rect 1835 -1222 2035 -1175
rect 2093 -1141 2293 -1125
rect 2093 -1175 2109 -1141
rect 2277 -1175 2293 -1141
rect 2093 -1222 2293 -1175
rect 2351 -1141 2551 -1125
rect 2351 -1175 2367 -1141
rect 2535 -1175 2551 -1141
rect 2351 -1222 2551 -1175
rect -2551 -1769 -2351 -1722
rect -2551 -1803 -2535 -1769
rect -2367 -1803 -2351 -1769
rect -2551 -1819 -2351 -1803
rect -2293 -1769 -2093 -1722
rect -2293 -1803 -2277 -1769
rect -2109 -1803 -2093 -1769
rect -2293 -1819 -2093 -1803
rect -2035 -1769 -1835 -1722
rect -2035 -1803 -2019 -1769
rect -1851 -1803 -1835 -1769
rect -2035 -1819 -1835 -1803
rect -1777 -1769 -1577 -1722
rect -1777 -1803 -1761 -1769
rect -1593 -1803 -1577 -1769
rect -1777 -1819 -1577 -1803
rect -1519 -1769 -1319 -1722
rect -1519 -1803 -1503 -1769
rect -1335 -1803 -1319 -1769
rect -1519 -1819 -1319 -1803
rect -1261 -1769 -1061 -1722
rect -1261 -1803 -1245 -1769
rect -1077 -1803 -1061 -1769
rect -1261 -1819 -1061 -1803
rect -1003 -1769 -803 -1722
rect -1003 -1803 -987 -1769
rect -819 -1803 -803 -1769
rect -1003 -1819 -803 -1803
rect -745 -1769 -545 -1722
rect -745 -1803 -729 -1769
rect -561 -1803 -545 -1769
rect -745 -1819 -545 -1803
rect -487 -1769 -287 -1722
rect -487 -1803 -471 -1769
rect -303 -1803 -287 -1769
rect -487 -1819 -287 -1803
rect -229 -1769 -29 -1722
rect -229 -1803 -213 -1769
rect -45 -1803 -29 -1769
rect -229 -1819 -29 -1803
rect 29 -1769 229 -1722
rect 29 -1803 45 -1769
rect 213 -1803 229 -1769
rect 29 -1819 229 -1803
rect 287 -1769 487 -1722
rect 287 -1803 303 -1769
rect 471 -1803 487 -1769
rect 287 -1819 487 -1803
rect 545 -1769 745 -1722
rect 545 -1803 561 -1769
rect 729 -1803 745 -1769
rect 545 -1819 745 -1803
rect 803 -1769 1003 -1722
rect 803 -1803 819 -1769
rect 987 -1803 1003 -1769
rect 803 -1819 1003 -1803
rect 1061 -1769 1261 -1722
rect 1061 -1803 1077 -1769
rect 1245 -1803 1261 -1769
rect 1061 -1819 1261 -1803
rect 1319 -1769 1519 -1722
rect 1319 -1803 1335 -1769
rect 1503 -1803 1519 -1769
rect 1319 -1819 1519 -1803
rect 1577 -1769 1777 -1722
rect 1577 -1803 1593 -1769
rect 1761 -1803 1777 -1769
rect 1577 -1819 1777 -1803
rect 1835 -1769 2035 -1722
rect 1835 -1803 1851 -1769
rect 2019 -1803 2035 -1769
rect 1835 -1819 2035 -1803
rect 2093 -1769 2293 -1722
rect 2093 -1803 2109 -1769
rect 2277 -1803 2293 -1769
rect 2093 -1819 2293 -1803
rect 2351 -1769 2551 -1722
rect 2351 -1803 2367 -1769
rect 2535 -1803 2551 -1769
rect 2351 -1819 2551 -1803
rect -2551 -1877 -2351 -1861
rect -2551 -1911 -2535 -1877
rect -2367 -1911 -2351 -1877
rect -2551 -1958 -2351 -1911
rect -2293 -1877 -2093 -1861
rect -2293 -1911 -2277 -1877
rect -2109 -1911 -2093 -1877
rect -2293 -1958 -2093 -1911
rect -2035 -1877 -1835 -1861
rect -2035 -1911 -2019 -1877
rect -1851 -1911 -1835 -1877
rect -2035 -1958 -1835 -1911
rect -1777 -1877 -1577 -1861
rect -1777 -1911 -1761 -1877
rect -1593 -1911 -1577 -1877
rect -1777 -1958 -1577 -1911
rect -1519 -1877 -1319 -1861
rect -1519 -1911 -1503 -1877
rect -1335 -1911 -1319 -1877
rect -1519 -1958 -1319 -1911
rect -1261 -1877 -1061 -1861
rect -1261 -1911 -1245 -1877
rect -1077 -1911 -1061 -1877
rect -1261 -1958 -1061 -1911
rect -1003 -1877 -803 -1861
rect -1003 -1911 -987 -1877
rect -819 -1911 -803 -1877
rect -1003 -1958 -803 -1911
rect -745 -1877 -545 -1861
rect -745 -1911 -729 -1877
rect -561 -1911 -545 -1877
rect -745 -1958 -545 -1911
rect -487 -1877 -287 -1861
rect -487 -1911 -471 -1877
rect -303 -1911 -287 -1877
rect -487 -1958 -287 -1911
rect -229 -1877 -29 -1861
rect -229 -1911 -213 -1877
rect -45 -1911 -29 -1877
rect -229 -1958 -29 -1911
rect 29 -1877 229 -1861
rect 29 -1911 45 -1877
rect 213 -1911 229 -1877
rect 29 -1958 229 -1911
rect 287 -1877 487 -1861
rect 287 -1911 303 -1877
rect 471 -1911 487 -1877
rect 287 -1958 487 -1911
rect 545 -1877 745 -1861
rect 545 -1911 561 -1877
rect 729 -1911 745 -1877
rect 545 -1958 745 -1911
rect 803 -1877 1003 -1861
rect 803 -1911 819 -1877
rect 987 -1911 1003 -1877
rect 803 -1958 1003 -1911
rect 1061 -1877 1261 -1861
rect 1061 -1911 1077 -1877
rect 1245 -1911 1261 -1877
rect 1061 -1958 1261 -1911
rect 1319 -1877 1519 -1861
rect 1319 -1911 1335 -1877
rect 1503 -1911 1519 -1877
rect 1319 -1958 1519 -1911
rect 1577 -1877 1777 -1861
rect 1577 -1911 1593 -1877
rect 1761 -1911 1777 -1877
rect 1577 -1958 1777 -1911
rect 1835 -1877 2035 -1861
rect 1835 -1911 1851 -1877
rect 2019 -1911 2035 -1877
rect 1835 -1958 2035 -1911
rect 2093 -1877 2293 -1861
rect 2093 -1911 2109 -1877
rect 2277 -1911 2293 -1877
rect 2093 -1958 2293 -1911
rect 2351 -1877 2551 -1861
rect 2351 -1911 2367 -1877
rect 2535 -1911 2551 -1877
rect 2351 -1958 2551 -1911
rect -2551 -2505 -2351 -2458
rect -2551 -2539 -2535 -2505
rect -2367 -2539 -2351 -2505
rect -2551 -2555 -2351 -2539
rect -2293 -2505 -2093 -2458
rect -2293 -2539 -2277 -2505
rect -2109 -2539 -2093 -2505
rect -2293 -2555 -2093 -2539
rect -2035 -2505 -1835 -2458
rect -2035 -2539 -2019 -2505
rect -1851 -2539 -1835 -2505
rect -2035 -2555 -1835 -2539
rect -1777 -2505 -1577 -2458
rect -1777 -2539 -1761 -2505
rect -1593 -2539 -1577 -2505
rect -1777 -2555 -1577 -2539
rect -1519 -2505 -1319 -2458
rect -1519 -2539 -1503 -2505
rect -1335 -2539 -1319 -2505
rect -1519 -2555 -1319 -2539
rect -1261 -2505 -1061 -2458
rect -1261 -2539 -1245 -2505
rect -1077 -2539 -1061 -2505
rect -1261 -2555 -1061 -2539
rect -1003 -2505 -803 -2458
rect -1003 -2539 -987 -2505
rect -819 -2539 -803 -2505
rect -1003 -2555 -803 -2539
rect -745 -2505 -545 -2458
rect -745 -2539 -729 -2505
rect -561 -2539 -545 -2505
rect -745 -2555 -545 -2539
rect -487 -2505 -287 -2458
rect -487 -2539 -471 -2505
rect -303 -2539 -287 -2505
rect -487 -2555 -287 -2539
rect -229 -2505 -29 -2458
rect -229 -2539 -213 -2505
rect -45 -2539 -29 -2505
rect -229 -2555 -29 -2539
rect 29 -2505 229 -2458
rect 29 -2539 45 -2505
rect 213 -2539 229 -2505
rect 29 -2555 229 -2539
rect 287 -2505 487 -2458
rect 287 -2539 303 -2505
rect 471 -2539 487 -2505
rect 287 -2555 487 -2539
rect 545 -2505 745 -2458
rect 545 -2539 561 -2505
rect 729 -2539 745 -2505
rect 545 -2555 745 -2539
rect 803 -2505 1003 -2458
rect 803 -2539 819 -2505
rect 987 -2539 1003 -2505
rect 803 -2555 1003 -2539
rect 1061 -2505 1261 -2458
rect 1061 -2539 1077 -2505
rect 1245 -2539 1261 -2505
rect 1061 -2555 1261 -2539
rect 1319 -2505 1519 -2458
rect 1319 -2539 1335 -2505
rect 1503 -2539 1519 -2505
rect 1319 -2555 1519 -2539
rect 1577 -2505 1777 -2458
rect 1577 -2539 1593 -2505
rect 1761 -2539 1777 -2505
rect 1577 -2555 1777 -2539
rect 1835 -2505 2035 -2458
rect 1835 -2539 1851 -2505
rect 2019 -2539 2035 -2505
rect 1835 -2555 2035 -2539
rect 2093 -2505 2293 -2458
rect 2093 -2539 2109 -2505
rect 2277 -2539 2293 -2505
rect 2093 -2555 2293 -2539
rect 2351 -2505 2551 -2458
rect 2351 -2539 2367 -2505
rect 2535 -2539 2551 -2505
rect 2351 -2555 2551 -2539
<< polycont >>
rect -2535 2505 -2367 2539
rect -2277 2505 -2109 2539
rect -2019 2505 -1851 2539
rect -1761 2505 -1593 2539
rect -1503 2505 -1335 2539
rect -1245 2505 -1077 2539
rect -987 2505 -819 2539
rect -729 2505 -561 2539
rect -471 2505 -303 2539
rect -213 2505 -45 2539
rect 45 2505 213 2539
rect 303 2505 471 2539
rect 561 2505 729 2539
rect 819 2505 987 2539
rect 1077 2505 1245 2539
rect 1335 2505 1503 2539
rect 1593 2505 1761 2539
rect 1851 2505 2019 2539
rect 2109 2505 2277 2539
rect 2367 2505 2535 2539
rect -2535 1877 -2367 1911
rect -2277 1877 -2109 1911
rect -2019 1877 -1851 1911
rect -1761 1877 -1593 1911
rect -1503 1877 -1335 1911
rect -1245 1877 -1077 1911
rect -987 1877 -819 1911
rect -729 1877 -561 1911
rect -471 1877 -303 1911
rect -213 1877 -45 1911
rect 45 1877 213 1911
rect 303 1877 471 1911
rect 561 1877 729 1911
rect 819 1877 987 1911
rect 1077 1877 1245 1911
rect 1335 1877 1503 1911
rect 1593 1877 1761 1911
rect 1851 1877 2019 1911
rect 2109 1877 2277 1911
rect 2367 1877 2535 1911
rect -2535 1769 -2367 1803
rect -2277 1769 -2109 1803
rect -2019 1769 -1851 1803
rect -1761 1769 -1593 1803
rect -1503 1769 -1335 1803
rect -1245 1769 -1077 1803
rect -987 1769 -819 1803
rect -729 1769 -561 1803
rect -471 1769 -303 1803
rect -213 1769 -45 1803
rect 45 1769 213 1803
rect 303 1769 471 1803
rect 561 1769 729 1803
rect 819 1769 987 1803
rect 1077 1769 1245 1803
rect 1335 1769 1503 1803
rect 1593 1769 1761 1803
rect 1851 1769 2019 1803
rect 2109 1769 2277 1803
rect 2367 1769 2535 1803
rect -2535 1141 -2367 1175
rect -2277 1141 -2109 1175
rect -2019 1141 -1851 1175
rect -1761 1141 -1593 1175
rect -1503 1141 -1335 1175
rect -1245 1141 -1077 1175
rect -987 1141 -819 1175
rect -729 1141 -561 1175
rect -471 1141 -303 1175
rect -213 1141 -45 1175
rect 45 1141 213 1175
rect 303 1141 471 1175
rect 561 1141 729 1175
rect 819 1141 987 1175
rect 1077 1141 1245 1175
rect 1335 1141 1503 1175
rect 1593 1141 1761 1175
rect 1851 1141 2019 1175
rect 2109 1141 2277 1175
rect 2367 1141 2535 1175
rect -2535 1033 -2367 1067
rect -2277 1033 -2109 1067
rect -2019 1033 -1851 1067
rect -1761 1033 -1593 1067
rect -1503 1033 -1335 1067
rect -1245 1033 -1077 1067
rect -987 1033 -819 1067
rect -729 1033 -561 1067
rect -471 1033 -303 1067
rect -213 1033 -45 1067
rect 45 1033 213 1067
rect 303 1033 471 1067
rect 561 1033 729 1067
rect 819 1033 987 1067
rect 1077 1033 1245 1067
rect 1335 1033 1503 1067
rect 1593 1033 1761 1067
rect 1851 1033 2019 1067
rect 2109 1033 2277 1067
rect 2367 1033 2535 1067
rect -2535 405 -2367 439
rect -2277 405 -2109 439
rect -2019 405 -1851 439
rect -1761 405 -1593 439
rect -1503 405 -1335 439
rect -1245 405 -1077 439
rect -987 405 -819 439
rect -729 405 -561 439
rect -471 405 -303 439
rect -213 405 -45 439
rect 45 405 213 439
rect 303 405 471 439
rect 561 405 729 439
rect 819 405 987 439
rect 1077 405 1245 439
rect 1335 405 1503 439
rect 1593 405 1761 439
rect 1851 405 2019 439
rect 2109 405 2277 439
rect 2367 405 2535 439
rect -2535 297 -2367 331
rect -2277 297 -2109 331
rect -2019 297 -1851 331
rect -1761 297 -1593 331
rect -1503 297 -1335 331
rect -1245 297 -1077 331
rect -987 297 -819 331
rect -729 297 -561 331
rect -471 297 -303 331
rect -213 297 -45 331
rect 45 297 213 331
rect 303 297 471 331
rect 561 297 729 331
rect 819 297 987 331
rect 1077 297 1245 331
rect 1335 297 1503 331
rect 1593 297 1761 331
rect 1851 297 2019 331
rect 2109 297 2277 331
rect 2367 297 2535 331
rect -2535 -331 -2367 -297
rect -2277 -331 -2109 -297
rect -2019 -331 -1851 -297
rect -1761 -331 -1593 -297
rect -1503 -331 -1335 -297
rect -1245 -331 -1077 -297
rect -987 -331 -819 -297
rect -729 -331 -561 -297
rect -471 -331 -303 -297
rect -213 -331 -45 -297
rect 45 -331 213 -297
rect 303 -331 471 -297
rect 561 -331 729 -297
rect 819 -331 987 -297
rect 1077 -331 1245 -297
rect 1335 -331 1503 -297
rect 1593 -331 1761 -297
rect 1851 -331 2019 -297
rect 2109 -331 2277 -297
rect 2367 -331 2535 -297
rect -2535 -439 -2367 -405
rect -2277 -439 -2109 -405
rect -2019 -439 -1851 -405
rect -1761 -439 -1593 -405
rect -1503 -439 -1335 -405
rect -1245 -439 -1077 -405
rect -987 -439 -819 -405
rect -729 -439 -561 -405
rect -471 -439 -303 -405
rect -213 -439 -45 -405
rect 45 -439 213 -405
rect 303 -439 471 -405
rect 561 -439 729 -405
rect 819 -439 987 -405
rect 1077 -439 1245 -405
rect 1335 -439 1503 -405
rect 1593 -439 1761 -405
rect 1851 -439 2019 -405
rect 2109 -439 2277 -405
rect 2367 -439 2535 -405
rect -2535 -1067 -2367 -1033
rect -2277 -1067 -2109 -1033
rect -2019 -1067 -1851 -1033
rect -1761 -1067 -1593 -1033
rect -1503 -1067 -1335 -1033
rect -1245 -1067 -1077 -1033
rect -987 -1067 -819 -1033
rect -729 -1067 -561 -1033
rect -471 -1067 -303 -1033
rect -213 -1067 -45 -1033
rect 45 -1067 213 -1033
rect 303 -1067 471 -1033
rect 561 -1067 729 -1033
rect 819 -1067 987 -1033
rect 1077 -1067 1245 -1033
rect 1335 -1067 1503 -1033
rect 1593 -1067 1761 -1033
rect 1851 -1067 2019 -1033
rect 2109 -1067 2277 -1033
rect 2367 -1067 2535 -1033
rect -2535 -1175 -2367 -1141
rect -2277 -1175 -2109 -1141
rect -2019 -1175 -1851 -1141
rect -1761 -1175 -1593 -1141
rect -1503 -1175 -1335 -1141
rect -1245 -1175 -1077 -1141
rect -987 -1175 -819 -1141
rect -729 -1175 -561 -1141
rect -471 -1175 -303 -1141
rect -213 -1175 -45 -1141
rect 45 -1175 213 -1141
rect 303 -1175 471 -1141
rect 561 -1175 729 -1141
rect 819 -1175 987 -1141
rect 1077 -1175 1245 -1141
rect 1335 -1175 1503 -1141
rect 1593 -1175 1761 -1141
rect 1851 -1175 2019 -1141
rect 2109 -1175 2277 -1141
rect 2367 -1175 2535 -1141
rect -2535 -1803 -2367 -1769
rect -2277 -1803 -2109 -1769
rect -2019 -1803 -1851 -1769
rect -1761 -1803 -1593 -1769
rect -1503 -1803 -1335 -1769
rect -1245 -1803 -1077 -1769
rect -987 -1803 -819 -1769
rect -729 -1803 -561 -1769
rect -471 -1803 -303 -1769
rect -213 -1803 -45 -1769
rect 45 -1803 213 -1769
rect 303 -1803 471 -1769
rect 561 -1803 729 -1769
rect 819 -1803 987 -1769
rect 1077 -1803 1245 -1769
rect 1335 -1803 1503 -1769
rect 1593 -1803 1761 -1769
rect 1851 -1803 2019 -1769
rect 2109 -1803 2277 -1769
rect 2367 -1803 2535 -1769
rect -2535 -1911 -2367 -1877
rect -2277 -1911 -2109 -1877
rect -2019 -1911 -1851 -1877
rect -1761 -1911 -1593 -1877
rect -1503 -1911 -1335 -1877
rect -1245 -1911 -1077 -1877
rect -987 -1911 -819 -1877
rect -729 -1911 -561 -1877
rect -471 -1911 -303 -1877
rect -213 -1911 -45 -1877
rect 45 -1911 213 -1877
rect 303 -1911 471 -1877
rect 561 -1911 729 -1877
rect 819 -1911 987 -1877
rect 1077 -1911 1245 -1877
rect 1335 -1911 1503 -1877
rect 1593 -1911 1761 -1877
rect 1851 -1911 2019 -1877
rect 2109 -1911 2277 -1877
rect 2367 -1911 2535 -1877
rect -2535 -2539 -2367 -2505
rect -2277 -2539 -2109 -2505
rect -2019 -2539 -1851 -2505
rect -1761 -2539 -1593 -2505
rect -1503 -2539 -1335 -2505
rect -1245 -2539 -1077 -2505
rect -987 -2539 -819 -2505
rect -729 -2539 -561 -2505
rect -471 -2539 -303 -2505
rect -213 -2539 -45 -2505
rect 45 -2539 213 -2505
rect 303 -2539 471 -2505
rect 561 -2539 729 -2505
rect 819 -2539 987 -2505
rect 1077 -2539 1245 -2505
rect 1335 -2539 1503 -2505
rect 1593 -2539 1761 -2505
rect 1851 -2539 2019 -2505
rect 2109 -2539 2277 -2505
rect 2367 -2539 2535 -2505
<< locali >>
rect -2711 2607 -2615 2641
rect 2615 2607 2711 2641
rect -2711 2545 -2677 2607
rect 2677 2545 2711 2607
rect -2551 2505 -2535 2539
rect -2367 2505 -2351 2539
rect -2293 2505 -2277 2539
rect -2109 2505 -2093 2539
rect -2035 2505 -2019 2539
rect -1851 2505 -1835 2539
rect -1777 2505 -1761 2539
rect -1593 2505 -1577 2539
rect -1519 2505 -1503 2539
rect -1335 2505 -1319 2539
rect -1261 2505 -1245 2539
rect -1077 2505 -1061 2539
rect -1003 2505 -987 2539
rect -819 2505 -803 2539
rect -745 2505 -729 2539
rect -561 2505 -545 2539
rect -487 2505 -471 2539
rect -303 2505 -287 2539
rect -229 2505 -213 2539
rect -45 2505 -29 2539
rect 29 2505 45 2539
rect 213 2505 229 2539
rect 287 2505 303 2539
rect 471 2505 487 2539
rect 545 2505 561 2539
rect 729 2505 745 2539
rect 803 2505 819 2539
rect 987 2505 1003 2539
rect 1061 2505 1077 2539
rect 1245 2505 1261 2539
rect 1319 2505 1335 2539
rect 1503 2505 1519 2539
rect 1577 2505 1593 2539
rect 1761 2505 1777 2539
rect 1835 2505 1851 2539
rect 2019 2505 2035 2539
rect 2093 2505 2109 2539
rect 2277 2505 2293 2539
rect 2351 2505 2367 2539
rect 2535 2505 2551 2539
rect -2597 2446 -2563 2462
rect -2597 1954 -2563 1970
rect -2339 2446 -2305 2462
rect -2339 1954 -2305 1970
rect -2081 2446 -2047 2462
rect -2081 1954 -2047 1970
rect -1823 2446 -1789 2462
rect -1823 1954 -1789 1970
rect -1565 2446 -1531 2462
rect -1565 1954 -1531 1970
rect -1307 2446 -1273 2462
rect -1307 1954 -1273 1970
rect -1049 2446 -1015 2462
rect -1049 1954 -1015 1970
rect -791 2446 -757 2462
rect -791 1954 -757 1970
rect -533 2446 -499 2462
rect -533 1954 -499 1970
rect -275 2446 -241 2462
rect -275 1954 -241 1970
rect -17 2446 17 2462
rect -17 1954 17 1970
rect 241 2446 275 2462
rect 241 1954 275 1970
rect 499 2446 533 2462
rect 499 1954 533 1970
rect 757 2446 791 2462
rect 757 1954 791 1970
rect 1015 2446 1049 2462
rect 1015 1954 1049 1970
rect 1273 2446 1307 2462
rect 1273 1954 1307 1970
rect 1531 2446 1565 2462
rect 1531 1954 1565 1970
rect 1789 2446 1823 2462
rect 1789 1954 1823 1970
rect 2047 2446 2081 2462
rect 2047 1954 2081 1970
rect 2305 2446 2339 2462
rect 2305 1954 2339 1970
rect 2563 2446 2597 2462
rect 2563 1954 2597 1970
rect -2551 1877 -2535 1911
rect -2367 1877 -2351 1911
rect -2293 1877 -2277 1911
rect -2109 1877 -2093 1911
rect -2035 1877 -2019 1911
rect -1851 1877 -1835 1911
rect -1777 1877 -1761 1911
rect -1593 1877 -1577 1911
rect -1519 1877 -1503 1911
rect -1335 1877 -1319 1911
rect -1261 1877 -1245 1911
rect -1077 1877 -1061 1911
rect -1003 1877 -987 1911
rect -819 1877 -803 1911
rect -745 1877 -729 1911
rect -561 1877 -545 1911
rect -487 1877 -471 1911
rect -303 1877 -287 1911
rect -229 1877 -213 1911
rect -45 1877 -29 1911
rect 29 1877 45 1911
rect 213 1877 229 1911
rect 287 1877 303 1911
rect 471 1877 487 1911
rect 545 1877 561 1911
rect 729 1877 745 1911
rect 803 1877 819 1911
rect 987 1877 1003 1911
rect 1061 1877 1077 1911
rect 1245 1877 1261 1911
rect 1319 1877 1335 1911
rect 1503 1877 1519 1911
rect 1577 1877 1593 1911
rect 1761 1877 1777 1911
rect 1835 1877 1851 1911
rect 2019 1877 2035 1911
rect 2093 1877 2109 1911
rect 2277 1877 2293 1911
rect 2351 1877 2367 1911
rect 2535 1877 2551 1911
rect -2551 1769 -2535 1803
rect -2367 1769 -2351 1803
rect -2293 1769 -2277 1803
rect -2109 1769 -2093 1803
rect -2035 1769 -2019 1803
rect -1851 1769 -1835 1803
rect -1777 1769 -1761 1803
rect -1593 1769 -1577 1803
rect -1519 1769 -1503 1803
rect -1335 1769 -1319 1803
rect -1261 1769 -1245 1803
rect -1077 1769 -1061 1803
rect -1003 1769 -987 1803
rect -819 1769 -803 1803
rect -745 1769 -729 1803
rect -561 1769 -545 1803
rect -487 1769 -471 1803
rect -303 1769 -287 1803
rect -229 1769 -213 1803
rect -45 1769 -29 1803
rect 29 1769 45 1803
rect 213 1769 229 1803
rect 287 1769 303 1803
rect 471 1769 487 1803
rect 545 1769 561 1803
rect 729 1769 745 1803
rect 803 1769 819 1803
rect 987 1769 1003 1803
rect 1061 1769 1077 1803
rect 1245 1769 1261 1803
rect 1319 1769 1335 1803
rect 1503 1769 1519 1803
rect 1577 1769 1593 1803
rect 1761 1769 1777 1803
rect 1835 1769 1851 1803
rect 2019 1769 2035 1803
rect 2093 1769 2109 1803
rect 2277 1769 2293 1803
rect 2351 1769 2367 1803
rect 2535 1769 2551 1803
rect -2597 1710 -2563 1726
rect -2597 1218 -2563 1234
rect -2339 1710 -2305 1726
rect -2339 1218 -2305 1234
rect -2081 1710 -2047 1726
rect -2081 1218 -2047 1234
rect -1823 1710 -1789 1726
rect -1823 1218 -1789 1234
rect -1565 1710 -1531 1726
rect -1565 1218 -1531 1234
rect -1307 1710 -1273 1726
rect -1307 1218 -1273 1234
rect -1049 1710 -1015 1726
rect -1049 1218 -1015 1234
rect -791 1710 -757 1726
rect -791 1218 -757 1234
rect -533 1710 -499 1726
rect -533 1218 -499 1234
rect -275 1710 -241 1726
rect -275 1218 -241 1234
rect -17 1710 17 1726
rect -17 1218 17 1234
rect 241 1710 275 1726
rect 241 1218 275 1234
rect 499 1710 533 1726
rect 499 1218 533 1234
rect 757 1710 791 1726
rect 757 1218 791 1234
rect 1015 1710 1049 1726
rect 1015 1218 1049 1234
rect 1273 1710 1307 1726
rect 1273 1218 1307 1234
rect 1531 1710 1565 1726
rect 1531 1218 1565 1234
rect 1789 1710 1823 1726
rect 1789 1218 1823 1234
rect 2047 1710 2081 1726
rect 2047 1218 2081 1234
rect 2305 1710 2339 1726
rect 2305 1218 2339 1234
rect 2563 1710 2597 1726
rect 2563 1218 2597 1234
rect -2551 1141 -2535 1175
rect -2367 1141 -2351 1175
rect -2293 1141 -2277 1175
rect -2109 1141 -2093 1175
rect -2035 1141 -2019 1175
rect -1851 1141 -1835 1175
rect -1777 1141 -1761 1175
rect -1593 1141 -1577 1175
rect -1519 1141 -1503 1175
rect -1335 1141 -1319 1175
rect -1261 1141 -1245 1175
rect -1077 1141 -1061 1175
rect -1003 1141 -987 1175
rect -819 1141 -803 1175
rect -745 1141 -729 1175
rect -561 1141 -545 1175
rect -487 1141 -471 1175
rect -303 1141 -287 1175
rect -229 1141 -213 1175
rect -45 1141 -29 1175
rect 29 1141 45 1175
rect 213 1141 229 1175
rect 287 1141 303 1175
rect 471 1141 487 1175
rect 545 1141 561 1175
rect 729 1141 745 1175
rect 803 1141 819 1175
rect 987 1141 1003 1175
rect 1061 1141 1077 1175
rect 1245 1141 1261 1175
rect 1319 1141 1335 1175
rect 1503 1141 1519 1175
rect 1577 1141 1593 1175
rect 1761 1141 1777 1175
rect 1835 1141 1851 1175
rect 2019 1141 2035 1175
rect 2093 1141 2109 1175
rect 2277 1141 2293 1175
rect 2351 1141 2367 1175
rect 2535 1141 2551 1175
rect -2551 1033 -2535 1067
rect -2367 1033 -2351 1067
rect -2293 1033 -2277 1067
rect -2109 1033 -2093 1067
rect -2035 1033 -2019 1067
rect -1851 1033 -1835 1067
rect -1777 1033 -1761 1067
rect -1593 1033 -1577 1067
rect -1519 1033 -1503 1067
rect -1335 1033 -1319 1067
rect -1261 1033 -1245 1067
rect -1077 1033 -1061 1067
rect -1003 1033 -987 1067
rect -819 1033 -803 1067
rect -745 1033 -729 1067
rect -561 1033 -545 1067
rect -487 1033 -471 1067
rect -303 1033 -287 1067
rect -229 1033 -213 1067
rect -45 1033 -29 1067
rect 29 1033 45 1067
rect 213 1033 229 1067
rect 287 1033 303 1067
rect 471 1033 487 1067
rect 545 1033 561 1067
rect 729 1033 745 1067
rect 803 1033 819 1067
rect 987 1033 1003 1067
rect 1061 1033 1077 1067
rect 1245 1033 1261 1067
rect 1319 1033 1335 1067
rect 1503 1033 1519 1067
rect 1577 1033 1593 1067
rect 1761 1033 1777 1067
rect 1835 1033 1851 1067
rect 2019 1033 2035 1067
rect 2093 1033 2109 1067
rect 2277 1033 2293 1067
rect 2351 1033 2367 1067
rect 2535 1033 2551 1067
rect -2597 974 -2563 990
rect -2597 482 -2563 498
rect -2339 974 -2305 990
rect -2339 482 -2305 498
rect -2081 974 -2047 990
rect -2081 482 -2047 498
rect -1823 974 -1789 990
rect -1823 482 -1789 498
rect -1565 974 -1531 990
rect -1565 482 -1531 498
rect -1307 974 -1273 990
rect -1307 482 -1273 498
rect -1049 974 -1015 990
rect -1049 482 -1015 498
rect -791 974 -757 990
rect -791 482 -757 498
rect -533 974 -499 990
rect -533 482 -499 498
rect -275 974 -241 990
rect -275 482 -241 498
rect -17 974 17 990
rect -17 482 17 498
rect 241 974 275 990
rect 241 482 275 498
rect 499 974 533 990
rect 499 482 533 498
rect 757 974 791 990
rect 757 482 791 498
rect 1015 974 1049 990
rect 1015 482 1049 498
rect 1273 974 1307 990
rect 1273 482 1307 498
rect 1531 974 1565 990
rect 1531 482 1565 498
rect 1789 974 1823 990
rect 1789 482 1823 498
rect 2047 974 2081 990
rect 2047 482 2081 498
rect 2305 974 2339 990
rect 2305 482 2339 498
rect 2563 974 2597 990
rect 2563 482 2597 498
rect -2551 405 -2535 439
rect -2367 405 -2351 439
rect -2293 405 -2277 439
rect -2109 405 -2093 439
rect -2035 405 -2019 439
rect -1851 405 -1835 439
rect -1777 405 -1761 439
rect -1593 405 -1577 439
rect -1519 405 -1503 439
rect -1335 405 -1319 439
rect -1261 405 -1245 439
rect -1077 405 -1061 439
rect -1003 405 -987 439
rect -819 405 -803 439
rect -745 405 -729 439
rect -561 405 -545 439
rect -487 405 -471 439
rect -303 405 -287 439
rect -229 405 -213 439
rect -45 405 -29 439
rect 29 405 45 439
rect 213 405 229 439
rect 287 405 303 439
rect 471 405 487 439
rect 545 405 561 439
rect 729 405 745 439
rect 803 405 819 439
rect 987 405 1003 439
rect 1061 405 1077 439
rect 1245 405 1261 439
rect 1319 405 1335 439
rect 1503 405 1519 439
rect 1577 405 1593 439
rect 1761 405 1777 439
rect 1835 405 1851 439
rect 2019 405 2035 439
rect 2093 405 2109 439
rect 2277 405 2293 439
rect 2351 405 2367 439
rect 2535 405 2551 439
rect -2551 297 -2535 331
rect -2367 297 -2351 331
rect -2293 297 -2277 331
rect -2109 297 -2093 331
rect -2035 297 -2019 331
rect -1851 297 -1835 331
rect -1777 297 -1761 331
rect -1593 297 -1577 331
rect -1519 297 -1503 331
rect -1335 297 -1319 331
rect -1261 297 -1245 331
rect -1077 297 -1061 331
rect -1003 297 -987 331
rect -819 297 -803 331
rect -745 297 -729 331
rect -561 297 -545 331
rect -487 297 -471 331
rect -303 297 -287 331
rect -229 297 -213 331
rect -45 297 -29 331
rect 29 297 45 331
rect 213 297 229 331
rect 287 297 303 331
rect 471 297 487 331
rect 545 297 561 331
rect 729 297 745 331
rect 803 297 819 331
rect 987 297 1003 331
rect 1061 297 1077 331
rect 1245 297 1261 331
rect 1319 297 1335 331
rect 1503 297 1519 331
rect 1577 297 1593 331
rect 1761 297 1777 331
rect 1835 297 1851 331
rect 2019 297 2035 331
rect 2093 297 2109 331
rect 2277 297 2293 331
rect 2351 297 2367 331
rect 2535 297 2551 331
rect -2597 238 -2563 254
rect -2597 -254 -2563 -238
rect -2339 238 -2305 254
rect -2339 -254 -2305 -238
rect -2081 238 -2047 254
rect -2081 -254 -2047 -238
rect -1823 238 -1789 254
rect -1823 -254 -1789 -238
rect -1565 238 -1531 254
rect -1565 -254 -1531 -238
rect -1307 238 -1273 254
rect -1307 -254 -1273 -238
rect -1049 238 -1015 254
rect -1049 -254 -1015 -238
rect -791 238 -757 254
rect -791 -254 -757 -238
rect -533 238 -499 254
rect -533 -254 -499 -238
rect -275 238 -241 254
rect -275 -254 -241 -238
rect -17 238 17 254
rect -17 -254 17 -238
rect 241 238 275 254
rect 241 -254 275 -238
rect 499 238 533 254
rect 499 -254 533 -238
rect 757 238 791 254
rect 757 -254 791 -238
rect 1015 238 1049 254
rect 1015 -254 1049 -238
rect 1273 238 1307 254
rect 1273 -254 1307 -238
rect 1531 238 1565 254
rect 1531 -254 1565 -238
rect 1789 238 1823 254
rect 1789 -254 1823 -238
rect 2047 238 2081 254
rect 2047 -254 2081 -238
rect 2305 238 2339 254
rect 2305 -254 2339 -238
rect 2563 238 2597 254
rect 2563 -254 2597 -238
rect -2551 -331 -2535 -297
rect -2367 -331 -2351 -297
rect -2293 -331 -2277 -297
rect -2109 -331 -2093 -297
rect -2035 -331 -2019 -297
rect -1851 -331 -1835 -297
rect -1777 -331 -1761 -297
rect -1593 -331 -1577 -297
rect -1519 -331 -1503 -297
rect -1335 -331 -1319 -297
rect -1261 -331 -1245 -297
rect -1077 -331 -1061 -297
rect -1003 -331 -987 -297
rect -819 -331 -803 -297
rect -745 -331 -729 -297
rect -561 -331 -545 -297
rect -487 -331 -471 -297
rect -303 -331 -287 -297
rect -229 -331 -213 -297
rect -45 -331 -29 -297
rect 29 -331 45 -297
rect 213 -331 229 -297
rect 287 -331 303 -297
rect 471 -331 487 -297
rect 545 -331 561 -297
rect 729 -331 745 -297
rect 803 -331 819 -297
rect 987 -331 1003 -297
rect 1061 -331 1077 -297
rect 1245 -331 1261 -297
rect 1319 -331 1335 -297
rect 1503 -331 1519 -297
rect 1577 -331 1593 -297
rect 1761 -331 1777 -297
rect 1835 -331 1851 -297
rect 2019 -331 2035 -297
rect 2093 -331 2109 -297
rect 2277 -331 2293 -297
rect 2351 -331 2367 -297
rect 2535 -331 2551 -297
rect -2551 -439 -2535 -405
rect -2367 -439 -2351 -405
rect -2293 -439 -2277 -405
rect -2109 -439 -2093 -405
rect -2035 -439 -2019 -405
rect -1851 -439 -1835 -405
rect -1777 -439 -1761 -405
rect -1593 -439 -1577 -405
rect -1519 -439 -1503 -405
rect -1335 -439 -1319 -405
rect -1261 -439 -1245 -405
rect -1077 -439 -1061 -405
rect -1003 -439 -987 -405
rect -819 -439 -803 -405
rect -745 -439 -729 -405
rect -561 -439 -545 -405
rect -487 -439 -471 -405
rect -303 -439 -287 -405
rect -229 -439 -213 -405
rect -45 -439 -29 -405
rect 29 -439 45 -405
rect 213 -439 229 -405
rect 287 -439 303 -405
rect 471 -439 487 -405
rect 545 -439 561 -405
rect 729 -439 745 -405
rect 803 -439 819 -405
rect 987 -439 1003 -405
rect 1061 -439 1077 -405
rect 1245 -439 1261 -405
rect 1319 -439 1335 -405
rect 1503 -439 1519 -405
rect 1577 -439 1593 -405
rect 1761 -439 1777 -405
rect 1835 -439 1851 -405
rect 2019 -439 2035 -405
rect 2093 -439 2109 -405
rect 2277 -439 2293 -405
rect 2351 -439 2367 -405
rect 2535 -439 2551 -405
rect -2597 -498 -2563 -482
rect -2597 -990 -2563 -974
rect -2339 -498 -2305 -482
rect -2339 -990 -2305 -974
rect -2081 -498 -2047 -482
rect -2081 -990 -2047 -974
rect -1823 -498 -1789 -482
rect -1823 -990 -1789 -974
rect -1565 -498 -1531 -482
rect -1565 -990 -1531 -974
rect -1307 -498 -1273 -482
rect -1307 -990 -1273 -974
rect -1049 -498 -1015 -482
rect -1049 -990 -1015 -974
rect -791 -498 -757 -482
rect -791 -990 -757 -974
rect -533 -498 -499 -482
rect -533 -990 -499 -974
rect -275 -498 -241 -482
rect -275 -990 -241 -974
rect -17 -498 17 -482
rect -17 -990 17 -974
rect 241 -498 275 -482
rect 241 -990 275 -974
rect 499 -498 533 -482
rect 499 -990 533 -974
rect 757 -498 791 -482
rect 757 -990 791 -974
rect 1015 -498 1049 -482
rect 1015 -990 1049 -974
rect 1273 -498 1307 -482
rect 1273 -990 1307 -974
rect 1531 -498 1565 -482
rect 1531 -990 1565 -974
rect 1789 -498 1823 -482
rect 1789 -990 1823 -974
rect 2047 -498 2081 -482
rect 2047 -990 2081 -974
rect 2305 -498 2339 -482
rect 2305 -990 2339 -974
rect 2563 -498 2597 -482
rect 2563 -990 2597 -974
rect -2551 -1067 -2535 -1033
rect -2367 -1067 -2351 -1033
rect -2293 -1067 -2277 -1033
rect -2109 -1067 -2093 -1033
rect -2035 -1067 -2019 -1033
rect -1851 -1067 -1835 -1033
rect -1777 -1067 -1761 -1033
rect -1593 -1067 -1577 -1033
rect -1519 -1067 -1503 -1033
rect -1335 -1067 -1319 -1033
rect -1261 -1067 -1245 -1033
rect -1077 -1067 -1061 -1033
rect -1003 -1067 -987 -1033
rect -819 -1067 -803 -1033
rect -745 -1067 -729 -1033
rect -561 -1067 -545 -1033
rect -487 -1067 -471 -1033
rect -303 -1067 -287 -1033
rect -229 -1067 -213 -1033
rect -45 -1067 -29 -1033
rect 29 -1067 45 -1033
rect 213 -1067 229 -1033
rect 287 -1067 303 -1033
rect 471 -1067 487 -1033
rect 545 -1067 561 -1033
rect 729 -1067 745 -1033
rect 803 -1067 819 -1033
rect 987 -1067 1003 -1033
rect 1061 -1067 1077 -1033
rect 1245 -1067 1261 -1033
rect 1319 -1067 1335 -1033
rect 1503 -1067 1519 -1033
rect 1577 -1067 1593 -1033
rect 1761 -1067 1777 -1033
rect 1835 -1067 1851 -1033
rect 2019 -1067 2035 -1033
rect 2093 -1067 2109 -1033
rect 2277 -1067 2293 -1033
rect 2351 -1067 2367 -1033
rect 2535 -1067 2551 -1033
rect -2551 -1175 -2535 -1141
rect -2367 -1175 -2351 -1141
rect -2293 -1175 -2277 -1141
rect -2109 -1175 -2093 -1141
rect -2035 -1175 -2019 -1141
rect -1851 -1175 -1835 -1141
rect -1777 -1175 -1761 -1141
rect -1593 -1175 -1577 -1141
rect -1519 -1175 -1503 -1141
rect -1335 -1175 -1319 -1141
rect -1261 -1175 -1245 -1141
rect -1077 -1175 -1061 -1141
rect -1003 -1175 -987 -1141
rect -819 -1175 -803 -1141
rect -745 -1175 -729 -1141
rect -561 -1175 -545 -1141
rect -487 -1175 -471 -1141
rect -303 -1175 -287 -1141
rect -229 -1175 -213 -1141
rect -45 -1175 -29 -1141
rect 29 -1175 45 -1141
rect 213 -1175 229 -1141
rect 287 -1175 303 -1141
rect 471 -1175 487 -1141
rect 545 -1175 561 -1141
rect 729 -1175 745 -1141
rect 803 -1175 819 -1141
rect 987 -1175 1003 -1141
rect 1061 -1175 1077 -1141
rect 1245 -1175 1261 -1141
rect 1319 -1175 1335 -1141
rect 1503 -1175 1519 -1141
rect 1577 -1175 1593 -1141
rect 1761 -1175 1777 -1141
rect 1835 -1175 1851 -1141
rect 2019 -1175 2035 -1141
rect 2093 -1175 2109 -1141
rect 2277 -1175 2293 -1141
rect 2351 -1175 2367 -1141
rect 2535 -1175 2551 -1141
rect -2597 -1234 -2563 -1218
rect -2597 -1726 -2563 -1710
rect -2339 -1234 -2305 -1218
rect -2339 -1726 -2305 -1710
rect -2081 -1234 -2047 -1218
rect -2081 -1726 -2047 -1710
rect -1823 -1234 -1789 -1218
rect -1823 -1726 -1789 -1710
rect -1565 -1234 -1531 -1218
rect -1565 -1726 -1531 -1710
rect -1307 -1234 -1273 -1218
rect -1307 -1726 -1273 -1710
rect -1049 -1234 -1015 -1218
rect -1049 -1726 -1015 -1710
rect -791 -1234 -757 -1218
rect -791 -1726 -757 -1710
rect -533 -1234 -499 -1218
rect -533 -1726 -499 -1710
rect -275 -1234 -241 -1218
rect -275 -1726 -241 -1710
rect -17 -1234 17 -1218
rect -17 -1726 17 -1710
rect 241 -1234 275 -1218
rect 241 -1726 275 -1710
rect 499 -1234 533 -1218
rect 499 -1726 533 -1710
rect 757 -1234 791 -1218
rect 757 -1726 791 -1710
rect 1015 -1234 1049 -1218
rect 1015 -1726 1049 -1710
rect 1273 -1234 1307 -1218
rect 1273 -1726 1307 -1710
rect 1531 -1234 1565 -1218
rect 1531 -1726 1565 -1710
rect 1789 -1234 1823 -1218
rect 1789 -1726 1823 -1710
rect 2047 -1234 2081 -1218
rect 2047 -1726 2081 -1710
rect 2305 -1234 2339 -1218
rect 2305 -1726 2339 -1710
rect 2563 -1234 2597 -1218
rect 2563 -1726 2597 -1710
rect -2551 -1803 -2535 -1769
rect -2367 -1803 -2351 -1769
rect -2293 -1803 -2277 -1769
rect -2109 -1803 -2093 -1769
rect -2035 -1803 -2019 -1769
rect -1851 -1803 -1835 -1769
rect -1777 -1803 -1761 -1769
rect -1593 -1803 -1577 -1769
rect -1519 -1803 -1503 -1769
rect -1335 -1803 -1319 -1769
rect -1261 -1803 -1245 -1769
rect -1077 -1803 -1061 -1769
rect -1003 -1803 -987 -1769
rect -819 -1803 -803 -1769
rect -745 -1803 -729 -1769
rect -561 -1803 -545 -1769
rect -487 -1803 -471 -1769
rect -303 -1803 -287 -1769
rect -229 -1803 -213 -1769
rect -45 -1803 -29 -1769
rect 29 -1803 45 -1769
rect 213 -1803 229 -1769
rect 287 -1803 303 -1769
rect 471 -1803 487 -1769
rect 545 -1803 561 -1769
rect 729 -1803 745 -1769
rect 803 -1803 819 -1769
rect 987 -1803 1003 -1769
rect 1061 -1803 1077 -1769
rect 1245 -1803 1261 -1769
rect 1319 -1803 1335 -1769
rect 1503 -1803 1519 -1769
rect 1577 -1803 1593 -1769
rect 1761 -1803 1777 -1769
rect 1835 -1803 1851 -1769
rect 2019 -1803 2035 -1769
rect 2093 -1803 2109 -1769
rect 2277 -1803 2293 -1769
rect 2351 -1803 2367 -1769
rect 2535 -1803 2551 -1769
rect -2551 -1911 -2535 -1877
rect -2367 -1911 -2351 -1877
rect -2293 -1911 -2277 -1877
rect -2109 -1911 -2093 -1877
rect -2035 -1911 -2019 -1877
rect -1851 -1911 -1835 -1877
rect -1777 -1911 -1761 -1877
rect -1593 -1911 -1577 -1877
rect -1519 -1911 -1503 -1877
rect -1335 -1911 -1319 -1877
rect -1261 -1911 -1245 -1877
rect -1077 -1911 -1061 -1877
rect -1003 -1911 -987 -1877
rect -819 -1911 -803 -1877
rect -745 -1911 -729 -1877
rect -561 -1911 -545 -1877
rect -487 -1911 -471 -1877
rect -303 -1911 -287 -1877
rect -229 -1911 -213 -1877
rect -45 -1911 -29 -1877
rect 29 -1911 45 -1877
rect 213 -1911 229 -1877
rect 287 -1911 303 -1877
rect 471 -1911 487 -1877
rect 545 -1911 561 -1877
rect 729 -1911 745 -1877
rect 803 -1911 819 -1877
rect 987 -1911 1003 -1877
rect 1061 -1911 1077 -1877
rect 1245 -1911 1261 -1877
rect 1319 -1911 1335 -1877
rect 1503 -1911 1519 -1877
rect 1577 -1911 1593 -1877
rect 1761 -1911 1777 -1877
rect 1835 -1911 1851 -1877
rect 2019 -1911 2035 -1877
rect 2093 -1911 2109 -1877
rect 2277 -1911 2293 -1877
rect 2351 -1911 2367 -1877
rect 2535 -1911 2551 -1877
rect -2597 -1970 -2563 -1954
rect -2597 -2462 -2563 -2446
rect -2339 -1970 -2305 -1954
rect -2339 -2462 -2305 -2446
rect -2081 -1970 -2047 -1954
rect -2081 -2462 -2047 -2446
rect -1823 -1970 -1789 -1954
rect -1823 -2462 -1789 -2446
rect -1565 -1970 -1531 -1954
rect -1565 -2462 -1531 -2446
rect -1307 -1970 -1273 -1954
rect -1307 -2462 -1273 -2446
rect -1049 -1970 -1015 -1954
rect -1049 -2462 -1015 -2446
rect -791 -1970 -757 -1954
rect -791 -2462 -757 -2446
rect -533 -1970 -499 -1954
rect -533 -2462 -499 -2446
rect -275 -1970 -241 -1954
rect -275 -2462 -241 -2446
rect -17 -1970 17 -1954
rect -17 -2462 17 -2446
rect 241 -1970 275 -1954
rect 241 -2462 275 -2446
rect 499 -1970 533 -1954
rect 499 -2462 533 -2446
rect 757 -1970 791 -1954
rect 757 -2462 791 -2446
rect 1015 -1970 1049 -1954
rect 1015 -2462 1049 -2446
rect 1273 -1970 1307 -1954
rect 1273 -2462 1307 -2446
rect 1531 -1970 1565 -1954
rect 1531 -2462 1565 -2446
rect 1789 -1970 1823 -1954
rect 1789 -2462 1823 -2446
rect 2047 -1970 2081 -1954
rect 2047 -2462 2081 -2446
rect 2305 -1970 2339 -1954
rect 2305 -2462 2339 -2446
rect 2563 -1970 2597 -1954
rect 2563 -2462 2597 -2446
rect -2551 -2539 -2535 -2505
rect -2367 -2539 -2351 -2505
rect -2293 -2539 -2277 -2505
rect -2109 -2539 -2093 -2505
rect -2035 -2539 -2019 -2505
rect -1851 -2539 -1835 -2505
rect -1777 -2539 -1761 -2505
rect -1593 -2539 -1577 -2505
rect -1519 -2539 -1503 -2505
rect -1335 -2539 -1319 -2505
rect -1261 -2539 -1245 -2505
rect -1077 -2539 -1061 -2505
rect -1003 -2539 -987 -2505
rect -819 -2539 -803 -2505
rect -745 -2539 -729 -2505
rect -561 -2539 -545 -2505
rect -487 -2539 -471 -2505
rect -303 -2539 -287 -2505
rect -229 -2539 -213 -2505
rect -45 -2539 -29 -2505
rect 29 -2539 45 -2505
rect 213 -2539 229 -2505
rect 287 -2539 303 -2505
rect 471 -2539 487 -2505
rect 545 -2539 561 -2505
rect 729 -2539 745 -2505
rect 803 -2539 819 -2505
rect 987 -2539 1003 -2505
rect 1061 -2539 1077 -2505
rect 1245 -2539 1261 -2505
rect 1319 -2539 1335 -2505
rect 1503 -2539 1519 -2505
rect 1577 -2539 1593 -2505
rect 1761 -2539 1777 -2505
rect 1835 -2539 1851 -2505
rect 2019 -2539 2035 -2505
rect 2093 -2539 2109 -2505
rect 2277 -2539 2293 -2505
rect 2351 -2539 2367 -2505
rect 2535 -2539 2551 -2505
rect -2711 -2607 -2677 -2545
rect 2677 -2607 2711 -2545
rect -2711 -2641 -2615 -2607
rect 2615 -2641 2711 -2607
<< viali >>
rect -2535 2505 -2367 2539
rect -2277 2505 -2109 2539
rect -2019 2505 -1851 2539
rect -1761 2505 -1593 2539
rect -1503 2505 -1335 2539
rect -1245 2505 -1077 2539
rect -987 2505 -819 2539
rect -729 2505 -561 2539
rect -471 2505 -303 2539
rect -213 2505 -45 2539
rect 45 2505 213 2539
rect 303 2505 471 2539
rect 561 2505 729 2539
rect 819 2505 987 2539
rect 1077 2505 1245 2539
rect 1335 2505 1503 2539
rect 1593 2505 1761 2539
rect 1851 2505 2019 2539
rect 2109 2505 2277 2539
rect 2367 2505 2535 2539
rect -2597 1970 -2563 2446
rect -2339 1970 -2305 2446
rect -2081 1970 -2047 2446
rect -1823 1970 -1789 2446
rect -1565 1970 -1531 2446
rect -1307 1970 -1273 2446
rect -1049 1970 -1015 2446
rect -791 1970 -757 2446
rect -533 1970 -499 2446
rect -275 1970 -241 2446
rect -17 1970 17 2446
rect 241 1970 275 2446
rect 499 1970 533 2446
rect 757 1970 791 2446
rect 1015 1970 1049 2446
rect 1273 1970 1307 2446
rect 1531 1970 1565 2446
rect 1789 1970 1823 2446
rect 2047 1970 2081 2446
rect 2305 1970 2339 2446
rect 2563 1970 2597 2446
rect -2535 1877 -2367 1911
rect -2277 1877 -2109 1911
rect -2019 1877 -1851 1911
rect -1761 1877 -1593 1911
rect -1503 1877 -1335 1911
rect -1245 1877 -1077 1911
rect -987 1877 -819 1911
rect -729 1877 -561 1911
rect -471 1877 -303 1911
rect -213 1877 -45 1911
rect 45 1877 213 1911
rect 303 1877 471 1911
rect 561 1877 729 1911
rect 819 1877 987 1911
rect 1077 1877 1245 1911
rect 1335 1877 1503 1911
rect 1593 1877 1761 1911
rect 1851 1877 2019 1911
rect 2109 1877 2277 1911
rect 2367 1877 2535 1911
rect -2535 1769 -2367 1803
rect -2277 1769 -2109 1803
rect -2019 1769 -1851 1803
rect -1761 1769 -1593 1803
rect -1503 1769 -1335 1803
rect -1245 1769 -1077 1803
rect -987 1769 -819 1803
rect -729 1769 -561 1803
rect -471 1769 -303 1803
rect -213 1769 -45 1803
rect 45 1769 213 1803
rect 303 1769 471 1803
rect 561 1769 729 1803
rect 819 1769 987 1803
rect 1077 1769 1245 1803
rect 1335 1769 1503 1803
rect 1593 1769 1761 1803
rect 1851 1769 2019 1803
rect 2109 1769 2277 1803
rect 2367 1769 2535 1803
rect -2597 1234 -2563 1710
rect -2339 1234 -2305 1710
rect -2081 1234 -2047 1710
rect -1823 1234 -1789 1710
rect -1565 1234 -1531 1710
rect -1307 1234 -1273 1710
rect -1049 1234 -1015 1710
rect -791 1234 -757 1710
rect -533 1234 -499 1710
rect -275 1234 -241 1710
rect -17 1234 17 1710
rect 241 1234 275 1710
rect 499 1234 533 1710
rect 757 1234 791 1710
rect 1015 1234 1049 1710
rect 1273 1234 1307 1710
rect 1531 1234 1565 1710
rect 1789 1234 1823 1710
rect 2047 1234 2081 1710
rect 2305 1234 2339 1710
rect 2563 1234 2597 1710
rect -2535 1141 -2367 1175
rect -2277 1141 -2109 1175
rect -2019 1141 -1851 1175
rect -1761 1141 -1593 1175
rect -1503 1141 -1335 1175
rect -1245 1141 -1077 1175
rect -987 1141 -819 1175
rect -729 1141 -561 1175
rect -471 1141 -303 1175
rect -213 1141 -45 1175
rect 45 1141 213 1175
rect 303 1141 471 1175
rect 561 1141 729 1175
rect 819 1141 987 1175
rect 1077 1141 1245 1175
rect 1335 1141 1503 1175
rect 1593 1141 1761 1175
rect 1851 1141 2019 1175
rect 2109 1141 2277 1175
rect 2367 1141 2535 1175
rect -2535 1033 -2367 1067
rect -2277 1033 -2109 1067
rect -2019 1033 -1851 1067
rect -1761 1033 -1593 1067
rect -1503 1033 -1335 1067
rect -1245 1033 -1077 1067
rect -987 1033 -819 1067
rect -729 1033 -561 1067
rect -471 1033 -303 1067
rect -213 1033 -45 1067
rect 45 1033 213 1067
rect 303 1033 471 1067
rect 561 1033 729 1067
rect 819 1033 987 1067
rect 1077 1033 1245 1067
rect 1335 1033 1503 1067
rect 1593 1033 1761 1067
rect 1851 1033 2019 1067
rect 2109 1033 2277 1067
rect 2367 1033 2535 1067
rect -2597 498 -2563 974
rect -2339 498 -2305 974
rect -2081 498 -2047 974
rect -1823 498 -1789 974
rect -1565 498 -1531 974
rect -1307 498 -1273 974
rect -1049 498 -1015 974
rect -791 498 -757 974
rect -533 498 -499 974
rect -275 498 -241 974
rect -17 498 17 974
rect 241 498 275 974
rect 499 498 533 974
rect 757 498 791 974
rect 1015 498 1049 974
rect 1273 498 1307 974
rect 1531 498 1565 974
rect 1789 498 1823 974
rect 2047 498 2081 974
rect 2305 498 2339 974
rect 2563 498 2597 974
rect -2535 405 -2367 439
rect -2277 405 -2109 439
rect -2019 405 -1851 439
rect -1761 405 -1593 439
rect -1503 405 -1335 439
rect -1245 405 -1077 439
rect -987 405 -819 439
rect -729 405 -561 439
rect -471 405 -303 439
rect -213 405 -45 439
rect 45 405 213 439
rect 303 405 471 439
rect 561 405 729 439
rect 819 405 987 439
rect 1077 405 1245 439
rect 1335 405 1503 439
rect 1593 405 1761 439
rect 1851 405 2019 439
rect 2109 405 2277 439
rect 2367 405 2535 439
rect -2535 297 -2367 331
rect -2277 297 -2109 331
rect -2019 297 -1851 331
rect -1761 297 -1593 331
rect -1503 297 -1335 331
rect -1245 297 -1077 331
rect -987 297 -819 331
rect -729 297 -561 331
rect -471 297 -303 331
rect -213 297 -45 331
rect 45 297 213 331
rect 303 297 471 331
rect 561 297 729 331
rect 819 297 987 331
rect 1077 297 1245 331
rect 1335 297 1503 331
rect 1593 297 1761 331
rect 1851 297 2019 331
rect 2109 297 2277 331
rect 2367 297 2535 331
rect -2597 -238 -2563 238
rect -2339 -238 -2305 238
rect -2081 -238 -2047 238
rect -1823 -238 -1789 238
rect -1565 -238 -1531 238
rect -1307 -238 -1273 238
rect -1049 -238 -1015 238
rect -791 -238 -757 238
rect -533 -238 -499 238
rect -275 -238 -241 238
rect -17 -238 17 238
rect 241 -238 275 238
rect 499 -238 533 238
rect 757 -238 791 238
rect 1015 -238 1049 238
rect 1273 -238 1307 238
rect 1531 -238 1565 238
rect 1789 -238 1823 238
rect 2047 -238 2081 238
rect 2305 -238 2339 238
rect 2563 -238 2597 238
rect -2535 -331 -2367 -297
rect -2277 -331 -2109 -297
rect -2019 -331 -1851 -297
rect -1761 -331 -1593 -297
rect -1503 -331 -1335 -297
rect -1245 -331 -1077 -297
rect -987 -331 -819 -297
rect -729 -331 -561 -297
rect -471 -331 -303 -297
rect -213 -331 -45 -297
rect 45 -331 213 -297
rect 303 -331 471 -297
rect 561 -331 729 -297
rect 819 -331 987 -297
rect 1077 -331 1245 -297
rect 1335 -331 1503 -297
rect 1593 -331 1761 -297
rect 1851 -331 2019 -297
rect 2109 -331 2277 -297
rect 2367 -331 2535 -297
rect -2535 -439 -2367 -405
rect -2277 -439 -2109 -405
rect -2019 -439 -1851 -405
rect -1761 -439 -1593 -405
rect -1503 -439 -1335 -405
rect -1245 -439 -1077 -405
rect -987 -439 -819 -405
rect -729 -439 -561 -405
rect -471 -439 -303 -405
rect -213 -439 -45 -405
rect 45 -439 213 -405
rect 303 -439 471 -405
rect 561 -439 729 -405
rect 819 -439 987 -405
rect 1077 -439 1245 -405
rect 1335 -439 1503 -405
rect 1593 -439 1761 -405
rect 1851 -439 2019 -405
rect 2109 -439 2277 -405
rect 2367 -439 2535 -405
rect -2597 -974 -2563 -498
rect -2339 -974 -2305 -498
rect -2081 -974 -2047 -498
rect -1823 -974 -1789 -498
rect -1565 -974 -1531 -498
rect -1307 -974 -1273 -498
rect -1049 -974 -1015 -498
rect -791 -974 -757 -498
rect -533 -974 -499 -498
rect -275 -974 -241 -498
rect -17 -974 17 -498
rect 241 -974 275 -498
rect 499 -974 533 -498
rect 757 -974 791 -498
rect 1015 -974 1049 -498
rect 1273 -974 1307 -498
rect 1531 -974 1565 -498
rect 1789 -974 1823 -498
rect 2047 -974 2081 -498
rect 2305 -974 2339 -498
rect 2563 -974 2597 -498
rect -2535 -1067 -2367 -1033
rect -2277 -1067 -2109 -1033
rect -2019 -1067 -1851 -1033
rect -1761 -1067 -1593 -1033
rect -1503 -1067 -1335 -1033
rect -1245 -1067 -1077 -1033
rect -987 -1067 -819 -1033
rect -729 -1067 -561 -1033
rect -471 -1067 -303 -1033
rect -213 -1067 -45 -1033
rect 45 -1067 213 -1033
rect 303 -1067 471 -1033
rect 561 -1067 729 -1033
rect 819 -1067 987 -1033
rect 1077 -1067 1245 -1033
rect 1335 -1067 1503 -1033
rect 1593 -1067 1761 -1033
rect 1851 -1067 2019 -1033
rect 2109 -1067 2277 -1033
rect 2367 -1067 2535 -1033
rect -2535 -1175 -2367 -1141
rect -2277 -1175 -2109 -1141
rect -2019 -1175 -1851 -1141
rect -1761 -1175 -1593 -1141
rect -1503 -1175 -1335 -1141
rect -1245 -1175 -1077 -1141
rect -987 -1175 -819 -1141
rect -729 -1175 -561 -1141
rect -471 -1175 -303 -1141
rect -213 -1175 -45 -1141
rect 45 -1175 213 -1141
rect 303 -1175 471 -1141
rect 561 -1175 729 -1141
rect 819 -1175 987 -1141
rect 1077 -1175 1245 -1141
rect 1335 -1175 1503 -1141
rect 1593 -1175 1761 -1141
rect 1851 -1175 2019 -1141
rect 2109 -1175 2277 -1141
rect 2367 -1175 2535 -1141
rect -2597 -1710 -2563 -1234
rect -2339 -1710 -2305 -1234
rect -2081 -1710 -2047 -1234
rect -1823 -1710 -1789 -1234
rect -1565 -1710 -1531 -1234
rect -1307 -1710 -1273 -1234
rect -1049 -1710 -1015 -1234
rect -791 -1710 -757 -1234
rect -533 -1710 -499 -1234
rect -275 -1710 -241 -1234
rect -17 -1710 17 -1234
rect 241 -1710 275 -1234
rect 499 -1710 533 -1234
rect 757 -1710 791 -1234
rect 1015 -1710 1049 -1234
rect 1273 -1710 1307 -1234
rect 1531 -1710 1565 -1234
rect 1789 -1710 1823 -1234
rect 2047 -1710 2081 -1234
rect 2305 -1710 2339 -1234
rect 2563 -1710 2597 -1234
rect -2535 -1803 -2367 -1769
rect -2277 -1803 -2109 -1769
rect -2019 -1803 -1851 -1769
rect -1761 -1803 -1593 -1769
rect -1503 -1803 -1335 -1769
rect -1245 -1803 -1077 -1769
rect -987 -1803 -819 -1769
rect -729 -1803 -561 -1769
rect -471 -1803 -303 -1769
rect -213 -1803 -45 -1769
rect 45 -1803 213 -1769
rect 303 -1803 471 -1769
rect 561 -1803 729 -1769
rect 819 -1803 987 -1769
rect 1077 -1803 1245 -1769
rect 1335 -1803 1503 -1769
rect 1593 -1803 1761 -1769
rect 1851 -1803 2019 -1769
rect 2109 -1803 2277 -1769
rect 2367 -1803 2535 -1769
rect -2535 -1911 -2367 -1877
rect -2277 -1911 -2109 -1877
rect -2019 -1911 -1851 -1877
rect -1761 -1911 -1593 -1877
rect -1503 -1911 -1335 -1877
rect -1245 -1911 -1077 -1877
rect -987 -1911 -819 -1877
rect -729 -1911 -561 -1877
rect -471 -1911 -303 -1877
rect -213 -1911 -45 -1877
rect 45 -1911 213 -1877
rect 303 -1911 471 -1877
rect 561 -1911 729 -1877
rect 819 -1911 987 -1877
rect 1077 -1911 1245 -1877
rect 1335 -1911 1503 -1877
rect 1593 -1911 1761 -1877
rect 1851 -1911 2019 -1877
rect 2109 -1911 2277 -1877
rect 2367 -1911 2535 -1877
rect -2597 -2446 -2563 -1970
rect -2339 -2446 -2305 -1970
rect -2081 -2446 -2047 -1970
rect -1823 -2446 -1789 -1970
rect -1565 -2446 -1531 -1970
rect -1307 -2446 -1273 -1970
rect -1049 -2446 -1015 -1970
rect -791 -2446 -757 -1970
rect -533 -2446 -499 -1970
rect -275 -2446 -241 -1970
rect -17 -2446 17 -1970
rect 241 -2446 275 -1970
rect 499 -2446 533 -1970
rect 757 -2446 791 -1970
rect 1015 -2446 1049 -1970
rect 1273 -2446 1307 -1970
rect 1531 -2446 1565 -1970
rect 1789 -2446 1823 -1970
rect 2047 -2446 2081 -1970
rect 2305 -2446 2339 -1970
rect 2563 -2446 2597 -1970
rect -2535 -2539 -2367 -2505
rect -2277 -2539 -2109 -2505
rect -2019 -2539 -1851 -2505
rect -1761 -2539 -1593 -2505
rect -1503 -2539 -1335 -2505
rect -1245 -2539 -1077 -2505
rect -987 -2539 -819 -2505
rect -729 -2539 -561 -2505
rect -471 -2539 -303 -2505
rect -213 -2539 -45 -2505
rect 45 -2539 213 -2505
rect 303 -2539 471 -2505
rect 561 -2539 729 -2505
rect 819 -2539 987 -2505
rect 1077 -2539 1245 -2505
rect 1335 -2539 1503 -2505
rect 1593 -2539 1761 -2505
rect 1851 -2539 2019 -2505
rect 2109 -2539 2277 -2505
rect 2367 -2539 2535 -2505
<< metal1 >>
rect -2547 2539 -2355 2545
rect -2547 2505 -2535 2539
rect -2367 2505 -2355 2539
rect -2547 2499 -2355 2505
rect -2289 2539 -2097 2545
rect -2289 2505 -2277 2539
rect -2109 2505 -2097 2539
rect -2289 2499 -2097 2505
rect -2031 2539 -1839 2545
rect -2031 2505 -2019 2539
rect -1851 2505 -1839 2539
rect -2031 2499 -1839 2505
rect -1773 2539 -1581 2545
rect -1773 2505 -1761 2539
rect -1593 2505 -1581 2539
rect -1773 2499 -1581 2505
rect -1515 2539 -1323 2545
rect -1515 2505 -1503 2539
rect -1335 2505 -1323 2539
rect -1515 2499 -1323 2505
rect -1257 2539 -1065 2545
rect -1257 2505 -1245 2539
rect -1077 2505 -1065 2539
rect -1257 2499 -1065 2505
rect -999 2539 -807 2545
rect -999 2505 -987 2539
rect -819 2505 -807 2539
rect -999 2499 -807 2505
rect -741 2539 -549 2545
rect -741 2505 -729 2539
rect -561 2505 -549 2539
rect -741 2499 -549 2505
rect -483 2539 -291 2545
rect -483 2505 -471 2539
rect -303 2505 -291 2539
rect -483 2499 -291 2505
rect -225 2539 -33 2545
rect -225 2505 -213 2539
rect -45 2505 -33 2539
rect -225 2499 -33 2505
rect 33 2539 225 2545
rect 33 2505 45 2539
rect 213 2505 225 2539
rect 33 2499 225 2505
rect 291 2539 483 2545
rect 291 2505 303 2539
rect 471 2505 483 2539
rect 291 2499 483 2505
rect 549 2539 741 2545
rect 549 2505 561 2539
rect 729 2505 741 2539
rect 549 2499 741 2505
rect 807 2539 999 2545
rect 807 2505 819 2539
rect 987 2505 999 2539
rect 807 2499 999 2505
rect 1065 2539 1257 2545
rect 1065 2505 1077 2539
rect 1245 2505 1257 2539
rect 1065 2499 1257 2505
rect 1323 2539 1515 2545
rect 1323 2505 1335 2539
rect 1503 2505 1515 2539
rect 1323 2499 1515 2505
rect 1581 2539 1773 2545
rect 1581 2505 1593 2539
rect 1761 2505 1773 2539
rect 1581 2499 1773 2505
rect 1839 2539 2031 2545
rect 1839 2505 1851 2539
rect 2019 2505 2031 2539
rect 1839 2499 2031 2505
rect 2097 2539 2289 2545
rect 2097 2505 2109 2539
rect 2277 2505 2289 2539
rect 2097 2499 2289 2505
rect 2355 2539 2547 2545
rect 2355 2505 2367 2539
rect 2535 2505 2547 2539
rect 2355 2499 2547 2505
rect -2603 2446 -2557 2458
rect -2603 1970 -2597 2446
rect -2563 1970 -2557 2446
rect -2603 1958 -2557 1970
rect -2345 2446 -2299 2458
rect -2345 1970 -2339 2446
rect -2305 1970 -2299 2446
rect -2345 1958 -2299 1970
rect -2087 2446 -2041 2458
rect -2087 1970 -2081 2446
rect -2047 1970 -2041 2446
rect -2087 1958 -2041 1970
rect -1829 2446 -1783 2458
rect -1829 1970 -1823 2446
rect -1789 1970 -1783 2446
rect -1829 1958 -1783 1970
rect -1571 2446 -1525 2458
rect -1571 1970 -1565 2446
rect -1531 1970 -1525 2446
rect -1571 1958 -1525 1970
rect -1313 2446 -1267 2458
rect -1313 1970 -1307 2446
rect -1273 1970 -1267 2446
rect -1313 1958 -1267 1970
rect -1055 2446 -1009 2458
rect -1055 1970 -1049 2446
rect -1015 1970 -1009 2446
rect -1055 1958 -1009 1970
rect -797 2446 -751 2458
rect -797 1970 -791 2446
rect -757 1970 -751 2446
rect -797 1958 -751 1970
rect -539 2446 -493 2458
rect -539 1970 -533 2446
rect -499 1970 -493 2446
rect -539 1958 -493 1970
rect -281 2446 -235 2458
rect -281 1970 -275 2446
rect -241 1970 -235 2446
rect -281 1958 -235 1970
rect -23 2446 23 2458
rect -23 1970 -17 2446
rect 17 1970 23 2446
rect -23 1958 23 1970
rect 235 2446 281 2458
rect 235 1970 241 2446
rect 275 1970 281 2446
rect 235 1958 281 1970
rect 493 2446 539 2458
rect 493 1970 499 2446
rect 533 1970 539 2446
rect 493 1958 539 1970
rect 751 2446 797 2458
rect 751 1970 757 2446
rect 791 1970 797 2446
rect 751 1958 797 1970
rect 1009 2446 1055 2458
rect 1009 1970 1015 2446
rect 1049 1970 1055 2446
rect 1009 1958 1055 1970
rect 1267 2446 1313 2458
rect 1267 1970 1273 2446
rect 1307 1970 1313 2446
rect 1267 1958 1313 1970
rect 1525 2446 1571 2458
rect 1525 1970 1531 2446
rect 1565 1970 1571 2446
rect 1525 1958 1571 1970
rect 1783 2446 1829 2458
rect 1783 1970 1789 2446
rect 1823 1970 1829 2446
rect 1783 1958 1829 1970
rect 2041 2446 2087 2458
rect 2041 1970 2047 2446
rect 2081 1970 2087 2446
rect 2041 1958 2087 1970
rect 2299 2446 2345 2458
rect 2299 1970 2305 2446
rect 2339 1970 2345 2446
rect 2299 1958 2345 1970
rect 2557 2446 2603 2458
rect 2557 1970 2563 2446
rect 2597 1970 2603 2446
rect 2557 1958 2603 1970
rect -2547 1911 -2355 1917
rect -2547 1877 -2535 1911
rect -2367 1877 -2355 1911
rect -2547 1871 -2355 1877
rect -2289 1911 -2097 1917
rect -2289 1877 -2277 1911
rect -2109 1877 -2097 1911
rect -2289 1871 -2097 1877
rect -2031 1911 -1839 1917
rect -2031 1877 -2019 1911
rect -1851 1877 -1839 1911
rect -2031 1871 -1839 1877
rect -1773 1911 -1581 1917
rect -1773 1877 -1761 1911
rect -1593 1877 -1581 1911
rect -1773 1871 -1581 1877
rect -1515 1911 -1323 1917
rect -1515 1877 -1503 1911
rect -1335 1877 -1323 1911
rect -1515 1871 -1323 1877
rect -1257 1911 -1065 1917
rect -1257 1877 -1245 1911
rect -1077 1877 -1065 1911
rect -1257 1871 -1065 1877
rect -999 1911 -807 1917
rect -999 1877 -987 1911
rect -819 1877 -807 1911
rect -999 1871 -807 1877
rect -741 1911 -549 1917
rect -741 1877 -729 1911
rect -561 1877 -549 1911
rect -741 1871 -549 1877
rect -483 1911 -291 1917
rect -483 1877 -471 1911
rect -303 1877 -291 1911
rect -483 1871 -291 1877
rect -225 1911 -33 1917
rect -225 1877 -213 1911
rect -45 1877 -33 1911
rect -225 1871 -33 1877
rect 33 1911 225 1917
rect 33 1877 45 1911
rect 213 1877 225 1911
rect 33 1871 225 1877
rect 291 1911 483 1917
rect 291 1877 303 1911
rect 471 1877 483 1911
rect 291 1871 483 1877
rect 549 1911 741 1917
rect 549 1877 561 1911
rect 729 1877 741 1911
rect 549 1871 741 1877
rect 807 1911 999 1917
rect 807 1877 819 1911
rect 987 1877 999 1911
rect 807 1871 999 1877
rect 1065 1911 1257 1917
rect 1065 1877 1077 1911
rect 1245 1877 1257 1911
rect 1065 1871 1257 1877
rect 1323 1911 1515 1917
rect 1323 1877 1335 1911
rect 1503 1877 1515 1911
rect 1323 1871 1515 1877
rect 1581 1911 1773 1917
rect 1581 1877 1593 1911
rect 1761 1877 1773 1911
rect 1581 1871 1773 1877
rect 1839 1911 2031 1917
rect 1839 1877 1851 1911
rect 2019 1877 2031 1911
rect 1839 1871 2031 1877
rect 2097 1911 2289 1917
rect 2097 1877 2109 1911
rect 2277 1877 2289 1911
rect 2097 1871 2289 1877
rect 2355 1911 2547 1917
rect 2355 1877 2367 1911
rect 2535 1877 2547 1911
rect 2355 1871 2547 1877
rect -2547 1803 -2355 1809
rect -2547 1769 -2535 1803
rect -2367 1769 -2355 1803
rect -2547 1763 -2355 1769
rect -2289 1803 -2097 1809
rect -2289 1769 -2277 1803
rect -2109 1769 -2097 1803
rect -2289 1763 -2097 1769
rect -2031 1803 -1839 1809
rect -2031 1769 -2019 1803
rect -1851 1769 -1839 1803
rect -2031 1763 -1839 1769
rect -1773 1803 -1581 1809
rect -1773 1769 -1761 1803
rect -1593 1769 -1581 1803
rect -1773 1763 -1581 1769
rect -1515 1803 -1323 1809
rect -1515 1769 -1503 1803
rect -1335 1769 -1323 1803
rect -1515 1763 -1323 1769
rect -1257 1803 -1065 1809
rect -1257 1769 -1245 1803
rect -1077 1769 -1065 1803
rect -1257 1763 -1065 1769
rect -999 1803 -807 1809
rect -999 1769 -987 1803
rect -819 1769 -807 1803
rect -999 1763 -807 1769
rect -741 1803 -549 1809
rect -741 1769 -729 1803
rect -561 1769 -549 1803
rect -741 1763 -549 1769
rect -483 1803 -291 1809
rect -483 1769 -471 1803
rect -303 1769 -291 1803
rect -483 1763 -291 1769
rect -225 1803 -33 1809
rect -225 1769 -213 1803
rect -45 1769 -33 1803
rect -225 1763 -33 1769
rect 33 1803 225 1809
rect 33 1769 45 1803
rect 213 1769 225 1803
rect 33 1763 225 1769
rect 291 1803 483 1809
rect 291 1769 303 1803
rect 471 1769 483 1803
rect 291 1763 483 1769
rect 549 1803 741 1809
rect 549 1769 561 1803
rect 729 1769 741 1803
rect 549 1763 741 1769
rect 807 1803 999 1809
rect 807 1769 819 1803
rect 987 1769 999 1803
rect 807 1763 999 1769
rect 1065 1803 1257 1809
rect 1065 1769 1077 1803
rect 1245 1769 1257 1803
rect 1065 1763 1257 1769
rect 1323 1803 1515 1809
rect 1323 1769 1335 1803
rect 1503 1769 1515 1803
rect 1323 1763 1515 1769
rect 1581 1803 1773 1809
rect 1581 1769 1593 1803
rect 1761 1769 1773 1803
rect 1581 1763 1773 1769
rect 1839 1803 2031 1809
rect 1839 1769 1851 1803
rect 2019 1769 2031 1803
rect 1839 1763 2031 1769
rect 2097 1803 2289 1809
rect 2097 1769 2109 1803
rect 2277 1769 2289 1803
rect 2097 1763 2289 1769
rect 2355 1803 2547 1809
rect 2355 1769 2367 1803
rect 2535 1769 2547 1803
rect 2355 1763 2547 1769
rect -2603 1710 -2557 1722
rect -2603 1234 -2597 1710
rect -2563 1234 -2557 1710
rect -2603 1222 -2557 1234
rect -2345 1710 -2299 1722
rect -2345 1234 -2339 1710
rect -2305 1234 -2299 1710
rect -2345 1222 -2299 1234
rect -2087 1710 -2041 1722
rect -2087 1234 -2081 1710
rect -2047 1234 -2041 1710
rect -2087 1222 -2041 1234
rect -1829 1710 -1783 1722
rect -1829 1234 -1823 1710
rect -1789 1234 -1783 1710
rect -1829 1222 -1783 1234
rect -1571 1710 -1525 1722
rect -1571 1234 -1565 1710
rect -1531 1234 -1525 1710
rect -1571 1222 -1525 1234
rect -1313 1710 -1267 1722
rect -1313 1234 -1307 1710
rect -1273 1234 -1267 1710
rect -1313 1222 -1267 1234
rect -1055 1710 -1009 1722
rect -1055 1234 -1049 1710
rect -1015 1234 -1009 1710
rect -1055 1222 -1009 1234
rect -797 1710 -751 1722
rect -797 1234 -791 1710
rect -757 1234 -751 1710
rect -797 1222 -751 1234
rect -539 1710 -493 1722
rect -539 1234 -533 1710
rect -499 1234 -493 1710
rect -539 1222 -493 1234
rect -281 1710 -235 1722
rect -281 1234 -275 1710
rect -241 1234 -235 1710
rect -281 1222 -235 1234
rect -23 1710 23 1722
rect -23 1234 -17 1710
rect 17 1234 23 1710
rect -23 1222 23 1234
rect 235 1710 281 1722
rect 235 1234 241 1710
rect 275 1234 281 1710
rect 235 1222 281 1234
rect 493 1710 539 1722
rect 493 1234 499 1710
rect 533 1234 539 1710
rect 493 1222 539 1234
rect 751 1710 797 1722
rect 751 1234 757 1710
rect 791 1234 797 1710
rect 751 1222 797 1234
rect 1009 1710 1055 1722
rect 1009 1234 1015 1710
rect 1049 1234 1055 1710
rect 1009 1222 1055 1234
rect 1267 1710 1313 1722
rect 1267 1234 1273 1710
rect 1307 1234 1313 1710
rect 1267 1222 1313 1234
rect 1525 1710 1571 1722
rect 1525 1234 1531 1710
rect 1565 1234 1571 1710
rect 1525 1222 1571 1234
rect 1783 1710 1829 1722
rect 1783 1234 1789 1710
rect 1823 1234 1829 1710
rect 1783 1222 1829 1234
rect 2041 1710 2087 1722
rect 2041 1234 2047 1710
rect 2081 1234 2087 1710
rect 2041 1222 2087 1234
rect 2299 1710 2345 1722
rect 2299 1234 2305 1710
rect 2339 1234 2345 1710
rect 2299 1222 2345 1234
rect 2557 1710 2603 1722
rect 2557 1234 2563 1710
rect 2597 1234 2603 1710
rect 2557 1222 2603 1234
rect -2547 1175 -2355 1181
rect -2547 1141 -2535 1175
rect -2367 1141 -2355 1175
rect -2547 1135 -2355 1141
rect -2289 1175 -2097 1181
rect -2289 1141 -2277 1175
rect -2109 1141 -2097 1175
rect -2289 1135 -2097 1141
rect -2031 1175 -1839 1181
rect -2031 1141 -2019 1175
rect -1851 1141 -1839 1175
rect -2031 1135 -1839 1141
rect -1773 1175 -1581 1181
rect -1773 1141 -1761 1175
rect -1593 1141 -1581 1175
rect -1773 1135 -1581 1141
rect -1515 1175 -1323 1181
rect -1515 1141 -1503 1175
rect -1335 1141 -1323 1175
rect -1515 1135 -1323 1141
rect -1257 1175 -1065 1181
rect -1257 1141 -1245 1175
rect -1077 1141 -1065 1175
rect -1257 1135 -1065 1141
rect -999 1175 -807 1181
rect -999 1141 -987 1175
rect -819 1141 -807 1175
rect -999 1135 -807 1141
rect -741 1175 -549 1181
rect -741 1141 -729 1175
rect -561 1141 -549 1175
rect -741 1135 -549 1141
rect -483 1175 -291 1181
rect -483 1141 -471 1175
rect -303 1141 -291 1175
rect -483 1135 -291 1141
rect -225 1175 -33 1181
rect -225 1141 -213 1175
rect -45 1141 -33 1175
rect -225 1135 -33 1141
rect 33 1175 225 1181
rect 33 1141 45 1175
rect 213 1141 225 1175
rect 33 1135 225 1141
rect 291 1175 483 1181
rect 291 1141 303 1175
rect 471 1141 483 1175
rect 291 1135 483 1141
rect 549 1175 741 1181
rect 549 1141 561 1175
rect 729 1141 741 1175
rect 549 1135 741 1141
rect 807 1175 999 1181
rect 807 1141 819 1175
rect 987 1141 999 1175
rect 807 1135 999 1141
rect 1065 1175 1257 1181
rect 1065 1141 1077 1175
rect 1245 1141 1257 1175
rect 1065 1135 1257 1141
rect 1323 1175 1515 1181
rect 1323 1141 1335 1175
rect 1503 1141 1515 1175
rect 1323 1135 1515 1141
rect 1581 1175 1773 1181
rect 1581 1141 1593 1175
rect 1761 1141 1773 1175
rect 1581 1135 1773 1141
rect 1839 1175 2031 1181
rect 1839 1141 1851 1175
rect 2019 1141 2031 1175
rect 1839 1135 2031 1141
rect 2097 1175 2289 1181
rect 2097 1141 2109 1175
rect 2277 1141 2289 1175
rect 2097 1135 2289 1141
rect 2355 1175 2547 1181
rect 2355 1141 2367 1175
rect 2535 1141 2547 1175
rect 2355 1135 2547 1141
rect -2547 1067 -2355 1073
rect -2547 1033 -2535 1067
rect -2367 1033 -2355 1067
rect -2547 1027 -2355 1033
rect -2289 1067 -2097 1073
rect -2289 1033 -2277 1067
rect -2109 1033 -2097 1067
rect -2289 1027 -2097 1033
rect -2031 1067 -1839 1073
rect -2031 1033 -2019 1067
rect -1851 1033 -1839 1067
rect -2031 1027 -1839 1033
rect -1773 1067 -1581 1073
rect -1773 1033 -1761 1067
rect -1593 1033 -1581 1067
rect -1773 1027 -1581 1033
rect -1515 1067 -1323 1073
rect -1515 1033 -1503 1067
rect -1335 1033 -1323 1067
rect -1515 1027 -1323 1033
rect -1257 1067 -1065 1073
rect -1257 1033 -1245 1067
rect -1077 1033 -1065 1067
rect -1257 1027 -1065 1033
rect -999 1067 -807 1073
rect -999 1033 -987 1067
rect -819 1033 -807 1067
rect -999 1027 -807 1033
rect -741 1067 -549 1073
rect -741 1033 -729 1067
rect -561 1033 -549 1067
rect -741 1027 -549 1033
rect -483 1067 -291 1073
rect -483 1033 -471 1067
rect -303 1033 -291 1067
rect -483 1027 -291 1033
rect -225 1067 -33 1073
rect -225 1033 -213 1067
rect -45 1033 -33 1067
rect -225 1027 -33 1033
rect 33 1067 225 1073
rect 33 1033 45 1067
rect 213 1033 225 1067
rect 33 1027 225 1033
rect 291 1067 483 1073
rect 291 1033 303 1067
rect 471 1033 483 1067
rect 291 1027 483 1033
rect 549 1067 741 1073
rect 549 1033 561 1067
rect 729 1033 741 1067
rect 549 1027 741 1033
rect 807 1067 999 1073
rect 807 1033 819 1067
rect 987 1033 999 1067
rect 807 1027 999 1033
rect 1065 1067 1257 1073
rect 1065 1033 1077 1067
rect 1245 1033 1257 1067
rect 1065 1027 1257 1033
rect 1323 1067 1515 1073
rect 1323 1033 1335 1067
rect 1503 1033 1515 1067
rect 1323 1027 1515 1033
rect 1581 1067 1773 1073
rect 1581 1033 1593 1067
rect 1761 1033 1773 1067
rect 1581 1027 1773 1033
rect 1839 1067 2031 1073
rect 1839 1033 1851 1067
rect 2019 1033 2031 1067
rect 1839 1027 2031 1033
rect 2097 1067 2289 1073
rect 2097 1033 2109 1067
rect 2277 1033 2289 1067
rect 2097 1027 2289 1033
rect 2355 1067 2547 1073
rect 2355 1033 2367 1067
rect 2535 1033 2547 1067
rect 2355 1027 2547 1033
rect -2603 974 -2557 986
rect -2603 498 -2597 974
rect -2563 498 -2557 974
rect -2603 486 -2557 498
rect -2345 974 -2299 986
rect -2345 498 -2339 974
rect -2305 498 -2299 974
rect -2345 486 -2299 498
rect -2087 974 -2041 986
rect -2087 498 -2081 974
rect -2047 498 -2041 974
rect -2087 486 -2041 498
rect -1829 974 -1783 986
rect -1829 498 -1823 974
rect -1789 498 -1783 974
rect -1829 486 -1783 498
rect -1571 974 -1525 986
rect -1571 498 -1565 974
rect -1531 498 -1525 974
rect -1571 486 -1525 498
rect -1313 974 -1267 986
rect -1313 498 -1307 974
rect -1273 498 -1267 974
rect -1313 486 -1267 498
rect -1055 974 -1009 986
rect -1055 498 -1049 974
rect -1015 498 -1009 974
rect -1055 486 -1009 498
rect -797 974 -751 986
rect -797 498 -791 974
rect -757 498 -751 974
rect -797 486 -751 498
rect -539 974 -493 986
rect -539 498 -533 974
rect -499 498 -493 974
rect -539 486 -493 498
rect -281 974 -235 986
rect -281 498 -275 974
rect -241 498 -235 974
rect -281 486 -235 498
rect -23 974 23 986
rect -23 498 -17 974
rect 17 498 23 974
rect -23 486 23 498
rect 235 974 281 986
rect 235 498 241 974
rect 275 498 281 974
rect 235 486 281 498
rect 493 974 539 986
rect 493 498 499 974
rect 533 498 539 974
rect 493 486 539 498
rect 751 974 797 986
rect 751 498 757 974
rect 791 498 797 974
rect 751 486 797 498
rect 1009 974 1055 986
rect 1009 498 1015 974
rect 1049 498 1055 974
rect 1009 486 1055 498
rect 1267 974 1313 986
rect 1267 498 1273 974
rect 1307 498 1313 974
rect 1267 486 1313 498
rect 1525 974 1571 986
rect 1525 498 1531 974
rect 1565 498 1571 974
rect 1525 486 1571 498
rect 1783 974 1829 986
rect 1783 498 1789 974
rect 1823 498 1829 974
rect 1783 486 1829 498
rect 2041 974 2087 986
rect 2041 498 2047 974
rect 2081 498 2087 974
rect 2041 486 2087 498
rect 2299 974 2345 986
rect 2299 498 2305 974
rect 2339 498 2345 974
rect 2299 486 2345 498
rect 2557 974 2603 986
rect 2557 498 2563 974
rect 2597 498 2603 974
rect 2557 486 2603 498
rect -2547 439 -2355 445
rect -2547 405 -2535 439
rect -2367 405 -2355 439
rect -2547 399 -2355 405
rect -2289 439 -2097 445
rect -2289 405 -2277 439
rect -2109 405 -2097 439
rect -2289 399 -2097 405
rect -2031 439 -1839 445
rect -2031 405 -2019 439
rect -1851 405 -1839 439
rect -2031 399 -1839 405
rect -1773 439 -1581 445
rect -1773 405 -1761 439
rect -1593 405 -1581 439
rect -1773 399 -1581 405
rect -1515 439 -1323 445
rect -1515 405 -1503 439
rect -1335 405 -1323 439
rect -1515 399 -1323 405
rect -1257 439 -1065 445
rect -1257 405 -1245 439
rect -1077 405 -1065 439
rect -1257 399 -1065 405
rect -999 439 -807 445
rect -999 405 -987 439
rect -819 405 -807 439
rect -999 399 -807 405
rect -741 439 -549 445
rect -741 405 -729 439
rect -561 405 -549 439
rect -741 399 -549 405
rect -483 439 -291 445
rect -483 405 -471 439
rect -303 405 -291 439
rect -483 399 -291 405
rect -225 439 -33 445
rect -225 405 -213 439
rect -45 405 -33 439
rect -225 399 -33 405
rect 33 439 225 445
rect 33 405 45 439
rect 213 405 225 439
rect 33 399 225 405
rect 291 439 483 445
rect 291 405 303 439
rect 471 405 483 439
rect 291 399 483 405
rect 549 439 741 445
rect 549 405 561 439
rect 729 405 741 439
rect 549 399 741 405
rect 807 439 999 445
rect 807 405 819 439
rect 987 405 999 439
rect 807 399 999 405
rect 1065 439 1257 445
rect 1065 405 1077 439
rect 1245 405 1257 439
rect 1065 399 1257 405
rect 1323 439 1515 445
rect 1323 405 1335 439
rect 1503 405 1515 439
rect 1323 399 1515 405
rect 1581 439 1773 445
rect 1581 405 1593 439
rect 1761 405 1773 439
rect 1581 399 1773 405
rect 1839 439 2031 445
rect 1839 405 1851 439
rect 2019 405 2031 439
rect 1839 399 2031 405
rect 2097 439 2289 445
rect 2097 405 2109 439
rect 2277 405 2289 439
rect 2097 399 2289 405
rect 2355 439 2547 445
rect 2355 405 2367 439
rect 2535 405 2547 439
rect 2355 399 2547 405
rect -2547 331 -2355 337
rect -2547 297 -2535 331
rect -2367 297 -2355 331
rect -2547 291 -2355 297
rect -2289 331 -2097 337
rect -2289 297 -2277 331
rect -2109 297 -2097 331
rect -2289 291 -2097 297
rect -2031 331 -1839 337
rect -2031 297 -2019 331
rect -1851 297 -1839 331
rect -2031 291 -1839 297
rect -1773 331 -1581 337
rect -1773 297 -1761 331
rect -1593 297 -1581 331
rect -1773 291 -1581 297
rect -1515 331 -1323 337
rect -1515 297 -1503 331
rect -1335 297 -1323 331
rect -1515 291 -1323 297
rect -1257 331 -1065 337
rect -1257 297 -1245 331
rect -1077 297 -1065 331
rect -1257 291 -1065 297
rect -999 331 -807 337
rect -999 297 -987 331
rect -819 297 -807 331
rect -999 291 -807 297
rect -741 331 -549 337
rect -741 297 -729 331
rect -561 297 -549 331
rect -741 291 -549 297
rect -483 331 -291 337
rect -483 297 -471 331
rect -303 297 -291 331
rect -483 291 -291 297
rect -225 331 -33 337
rect -225 297 -213 331
rect -45 297 -33 331
rect -225 291 -33 297
rect 33 331 225 337
rect 33 297 45 331
rect 213 297 225 331
rect 33 291 225 297
rect 291 331 483 337
rect 291 297 303 331
rect 471 297 483 331
rect 291 291 483 297
rect 549 331 741 337
rect 549 297 561 331
rect 729 297 741 331
rect 549 291 741 297
rect 807 331 999 337
rect 807 297 819 331
rect 987 297 999 331
rect 807 291 999 297
rect 1065 331 1257 337
rect 1065 297 1077 331
rect 1245 297 1257 331
rect 1065 291 1257 297
rect 1323 331 1515 337
rect 1323 297 1335 331
rect 1503 297 1515 331
rect 1323 291 1515 297
rect 1581 331 1773 337
rect 1581 297 1593 331
rect 1761 297 1773 331
rect 1581 291 1773 297
rect 1839 331 2031 337
rect 1839 297 1851 331
rect 2019 297 2031 331
rect 1839 291 2031 297
rect 2097 331 2289 337
rect 2097 297 2109 331
rect 2277 297 2289 331
rect 2097 291 2289 297
rect 2355 331 2547 337
rect 2355 297 2367 331
rect 2535 297 2547 331
rect 2355 291 2547 297
rect -2603 238 -2557 250
rect -2603 -238 -2597 238
rect -2563 -238 -2557 238
rect -2603 -250 -2557 -238
rect -2345 238 -2299 250
rect -2345 -238 -2339 238
rect -2305 -238 -2299 238
rect -2345 -250 -2299 -238
rect -2087 238 -2041 250
rect -2087 -238 -2081 238
rect -2047 -238 -2041 238
rect -2087 -250 -2041 -238
rect -1829 238 -1783 250
rect -1829 -238 -1823 238
rect -1789 -238 -1783 238
rect -1829 -250 -1783 -238
rect -1571 238 -1525 250
rect -1571 -238 -1565 238
rect -1531 -238 -1525 238
rect -1571 -250 -1525 -238
rect -1313 238 -1267 250
rect -1313 -238 -1307 238
rect -1273 -238 -1267 238
rect -1313 -250 -1267 -238
rect -1055 238 -1009 250
rect -1055 -238 -1049 238
rect -1015 -238 -1009 238
rect -1055 -250 -1009 -238
rect -797 238 -751 250
rect -797 -238 -791 238
rect -757 -238 -751 238
rect -797 -250 -751 -238
rect -539 238 -493 250
rect -539 -238 -533 238
rect -499 -238 -493 238
rect -539 -250 -493 -238
rect -281 238 -235 250
rect -281 -238 -275 238
rect -241 -238 -235 238
rect -281 -250 -235 -238
rect -23 238 23 250
rect -23 -238 -17 238
rect 17 -238 23 238
rect -23 -250 23 -238
rect 235 238 281 250
rect 235 -238 241 238
rect 275 -238 281 238
rect 235 -250 281 -238
rect 493 238 539 250
rect 493 -238 499 238
rect 533 -238 539 238
rect 493 -250 539 -238
rect 751 238 797 250
rect 751 -238 757 238
rect 791 -238 797 238
rect 751 -250 797 -238
rect 1009 238 1055 250
rect 1009 -238 1015 238
rect 1049 -238 1055 238
rect 1009 -250 1055 -238
rect 1267 238 1313 250
rect 1267 -238 1273 238
rect 1307 -238 1313 238
rect 1267 -250 1313 -238
rect 1525 238 1571 250
rect 1525 -238 1531 238
rect 1565 -238 1571 238
rect 1525 -250 1571 -238
rect 1783 238 1829 250
rect 1783 -238 1789 238
rect 1823 -238 1829 238
rect 1783 -250 1829 -238
rect 2041 238 2087 250
rect 2041 -238 2047 238
rect 2081 -238 2087 238
rect 2041 -250 2087 -238
rect 2299 238 2345 250
rect 2299 -238 2305 238
rect 2339 -238 2345 238
rect 2299 -250 2345 -238
rect 2557 238 2603 250
rect 2557 -238 2563 238
rect 2597 -238 2603 238
rect 2557 -250 2603 -238
rect -2547 -297 -2355 -291
rect -2547 -331 -2535 -297
rect -2367 -331 -2355 -297
rect -2547 -337 -2355 -331
rect -2289 -297 -2097 -291
rect -2289 -331 -2277 -297
rect -2109 -331 -2097 -297
rect -2289 -337 -2097 -331
rect -2031 -297 -1839 -291
rect -2031 -331 -2019 -297
rect -1851 -331 -1839 -297
rect -2031 -337 -1839 -331
rect -1773 -297 -1581 -291
rect -1773 -331 -1761 -297
rect -1593 -331 -1581 -297
rect -1773 -337 -1581 -331
rect -1515 -297 -1323 -291
rect -1515 -331 -1503 -297
rect -1335 -331 -1323 -297
rect -1515 -337 -1323 -331
rect -1257 -297 -1065 -291
rect -1257 -331 -1245 -297
rect -1077 -331 -1065 -297
rect -1257 -337 -1065 -331
rect -999 -297 -807 -291
rect -999 -331 -987 -297
rect -819 -331 -807 -297
rect -999 -337 -807 -331
rect -741 -297 -549 -291
rect -741 -331 -729 -297
rect -561 -331 -549 -297
rect -741 -337 -549 -331
rect -483 -297 -291 -291
rect -483 -331 -471 -297
rect -303 -331 -291 -297
rect -483 -337 -291 -331
rect -225 -297 -33 -291
rect -225 -331 -213 -297
rect -45 -331 -33 -297
rect -225 -337 -33 -331
rect 33 -297 225 -291
rect 33 -331 45 -297
rect 213 -331 225 -297
rect 33 -337 225 -331
rect 291 -297 483 -291
rect 291 -331 303 -297
rect 471 -331 483 -297
rect 291 -337 483 -331
rect 549 -297 741 -291
rect 549 -331 561 -297
rect 729 -331 741 -297
rect 549 -337 741 -331
rect 807 -297 999 -291
rect 807 -331 819 -297
rect 987 -331 999 -297
rect 807 -337 999 -331
rect 1065 -297 1257 -291
rect 1065 -331 1077 -297
rect 1245 -331 1257 -297
rect 1065 -337 1257 -331
rect 1323 -297 1515 -291
rect 1323 -331 1335 -297
rect 1503 -331 1515 -297
rect 1323 -337 1515 -331
rect 1581 -297 1773 -291
rect 1581 -331 1593 -297
rect 1761 -331 1773 -297
rect 1581 -337 1773 -331
rect 1839 -297 2031 -291
rect 1839 -331 1851 -297
rect 2019 -331 2031 -297
rect 1839 -337 2031 -331
rect 2097 -297 2289 -291
rect 2097 -331 2109 -297
rect 2277 -331 2289 -297
rect 2097 -337 2289 -331
rect 2355 -297 2547 -291
rect 2355 -331 2367 -297
rect 2535 -331 2547 -297
rect 2355 -337 2547 -331
rect -2547 -405 -2355 -399
rect -2547 -439 -2535 -405
rect -2367 -439 -2355 -405
rect -2547 -445 -2355 -439
rect -2289 -405 -2097 -399
rect -2289 -439 -2277 -405
rect -2109 -439 -2097 -405
rect -2289 -445 -2097 -439
rect -2031 -405 -1839 -399
rect -2031 -439 -2019 -405
rect -1851 -439 -1839 -405
rect -2031 -445 -1839 -439
rect -1773 -405 -1581 -399
rect -1773 -439 -1761 -405
rect -1593 -439 -1581 -405
rect -1773 -445 -1581 -439
rect -1515 -405 -1323 -399
rect -1515 -439 -1503 -405
rect -1335 -439 -1323 -405
rect -1515 -445 -1323 -439
rect -1257 -405 -1065 -399
rect -1257 -439 -1245 -405
rect -1077 -439 -1065 -405
rect -1257 -445 -1065 -439
rect -999 -405 -807 -399
rect -999 -439 -987 -405
rect -819 -439 -807 -405
rect -999 -445 -807 -439
rect -741 -405 -549 -399
rect -741 -439 -729 -405
rect -561 -439 -549 -405
rect -741 -445 -549 -439
rect -483 -405 -291 -399
rect -483 -439 -471 -405
rect -303 -439 -291 -405
rect -483 -445 -291 -439
rect -225 -405 -33 -399
rect -225 -439 -213 -405
rect -45 -439 -33 -405
rect -225 -445 -33 -439
rect 33 -405 225 -399
rect 33 -439 45 -405
rect 213 -439 225 -405
rect 33 -445 225 -439
rect 291 -405 483 -399
rect 291 -439 303 -405
rect 471 -439 483 -405
rect 291 -445 483 -439
rect 549 -405 741 -399
rect 549 -439 561 -405
rect 729 -439 741 -405
rect 549 -445 741 -439
rect 807 -405 999 -399
rect 807 -439 819 -405
rect 987 -439 999 -405
rect 807 -445 999 -439
rect 1065 -405 1257 -399
rect 1065 -439 1077 -405
rect 1245 -439 1257 -405
rect 1065 -445 1257 -439
rect 1323 -405 1515 -399
rect 1323 -439 1335 -405
rect 1503 -439 1515 -405
rect 1323 -445 1515 -439
rect 1581 -405 1773 -399
rect 1581 -439 1593 -405
rect 1761 -439 1773 -405
rect 1581 -445 1773 -439
rect 1839 -405 2031 -399
rect 1839 -439 1851 -405
rect 2019 -439 2031 -405
rect 1839 -445 2031 -439
rect 2097 -405 2289 -399
rect 2097 -439 2109 -405
rect 2277 -439 2289 -405
rect 2097 -445 2289 -439
rect 2355 -405 2547 -399
rect 2355 -439 2367 -405
rect 2535 -439 2547 -405
rect 2355 -445 2547 -439
rect -2603 -498 -2557 -486
rect -2603 -974 -2597 -498
rect -2563 -974 -2557 -498
rect -2603 -986 -2557 -974
rect -2345 -498 -2299 -486
rect -2345 -974 -2339 -498
rect -2305 -974 -2299 -498
rect -2345 -986 -2299 -974
rect -2087 -498 -2041 -486
rect -2087 -974 -2081 -498
rect -2047 -974 -2041 -498
rect -2087 -986 -2041 -974
rect -1829 -498 -1783 -486
rect -1829 -974 -1823 -498
rect -1789 -974 -1783 -498
rect -1829 -986 -1783 -974
rect -1571 -498 -1525 -486
rect -1571 -974 -1565 -498
rect -1531 -974 -1525 -498
rect -1571 -986 -1525 -974
rect -1313 -498 -1267 -486
rect -1313 -974 -1307 -498
rect -1273 -974 -1267 -498
rect -1313 -986 -1267 -974
rect -1055 -498 -1009 -486
rect -1055 -974 -1049 -498
rect -1015 -974 -1009 -498
rect -1055 -986 -1009 -974
rect -797 -498 -751 -486
rect -797 -974 -791 -498
rect -757 -974 -751 -498
rect -797 -986 -751 -974
rect -539 -498 -493 -486
rect -539 -974 -533 -498
rect -499 -974 -493 -498
rect -539 -986 -493 -974
rect -281 -498 -235 -486
rect -281 -974 -275 -498
rect -241 -974 -235 -498
rect -281 -986 -235 -974
rect -23 -498 23 -486
rect -23 -974 -17 -498
rect 17 -974 23 -498
rect -23 -986 23 -974
rect 235 -498 281 -486
rect 235 -974 241 -498
rect 275 -974 281 -498
rect 235 -986 281 -974
rect 493 -498 539 -486
rect 493 -974 499 -498
rect 533 -974 539 -498
rect 493 -986 539 -974
rect 751 -498 797 -486
rect 751 -974 757 -498
rect 791 -974 797 -498
rect 751 -986 797 -974
rect 1009 -498 1055 -486
rect 1009 -974 1015 -498
rect 1049 -974 1055 -498
rect 1009 -986 1055 -974
rect 1267 -498 1313 -486
rect 1267 -974 1273 -498
rect 1307 -974 1313 -498
rect 1267 -986 1313 -974
rect 1525 -498 1571 -486
rect 1525 -974 1531 -498
rect 1565 -974 1571 -498
rect 1525 -986 1571 -974
rect 1783 -498 1829 -486
rect 1783 -974 1789 -498
rect 1823 -974 1829 -498
rect 1783 -986 1829 -974
rect 2041 -498 2087 -486
rect 2041 -974 2047 -498
rect 2081 -974 2087 -498
rect 2041 -986 2087 -974
rect 2299 -498 2345 -486
rect 2299 -974 2305 -498
rect 2339 -974 2345 -498
rect 2299 -986 2345 -974
rect 2557 -498 2603 -486
rect 2557 -974 2563 -498
rect 2597 -974 2603 -498
rect 2557 -986 2603 -974
rect -2547 -1033 -2355 -1027
rect -2547 -1067 -2535 -1033
rect -2367 -1067 -2355 -1033
rect -2547 -1073 -2355 -1067
rect -2289 -1033 -2097 -1027
rect -2289 -1067 -2277 -1033
rect -2109 -1067 -2097 -1033
rect -2289 -1073 -2097 -1067
rect -2031 -1033 -1839 -1027
rect -2031 -1067 -2019 -1033
rect -1851 -1067 -1839 -1033
rect -2031 -1073 -1839 -1067
rect -1773 -1033 -1581 -1027
rect -1773 -1067 -1761 -1033
rect -1593 -1067 -1581 -1033
rect -1773 -1073 -1581 -1067
rect -1515 -1033 -1323 -1027
rect -1515 -1067 -1503 -1033
rect -1335 -1067 -1323 -1033
rect -1515 -1073 -1323 -1067
rect -1257 -1033 -1065 -1027
rect -1257 -1067 -1245 -1033
rect -1077 -1067 -1065 -1033
rect -1257 -1073 -1065 -1067
rect -999 -1033 -807 -1027
rect -999 -1067 -987 -1033
rect -819 -1067 -807 -1033
rect -999 -1073 -807 -1067
rect -741 -1033 -549 -1027
rect -741 -1067 -729 -1033
rect -561 -1067 -549 -1033
rect -741 -1073 -549 -1067
rect -483 -1033 -291 -1027
rect -483 -1067 -471 -1033
rect -303 -1067 -291 -1033
rect -483 -1073 -291 -1067
rect -225 -1033 -33 -1027
rect -225 -1067 -213 -1033
rect -45 -1067 -33 -1033
rect -225 -1073 -33 -1067
rect 33 -1033 225 -1027
rect 33 -1067 45 -1033
rect 213 -1067 225 -1033
rect 33 -1073 225 -1067
rect 291 -1033 483 -1027
rect 291 -1067 303 -1033
rect 471 -1067 483 -1033
rect 291 -1073 483 -1067
rect 549 -1033 741 -1027
rect 549 -1067 561 -1033
rect 729 -1067 741 -1033
rect 549 -1073 741 -1067
rect 807 -1033 999 -1027
rect 807 -1067 819 -1033
rect 987 -1067 999 -1033
rect 807 -1073 999 -1067
rect 1065 -1033 1257 -1027
rect 1065 -1067 1077 -1033
rect 1245 -1067 1257 -1033
rect 1065 -1073 1257 -1067
rect 1323 -1033 1515 -1027
rect 1323 -1067 1335 -1033
rect 1503 -1067 1515 -1033
rect 1323 -1073 1515 -1067
rect 1581 -1033 1773 -1027
rect 1581 -1067 1593 -1033
rect 1761 -1067 1773 -1033
rect 1581 -1073 1773 -1067
rect 1839 -1033 2031 -1027
rect 1839 -1067 1851 -1033
rect 2019 -1067 2031 -1033
rect 1839 -1073 2031 -1067
rect 2097 -1033 2289 -1027
rect 2097 -1067 2109 -1033
rect 2277 -1067 2289 -1033
rect 2097 -1073 2289 -1067
rect 2355 -1033 2547 -1027
rect 2355 -1067 2367 -1033
rect 2535 -1067 2547 -1033
rect 2355 -1073 2547 -1067
rect -2547 -1141 -2355 -1135
rect -2547 -1175 -2535 -1141
rect -2367 -1175 -2355 -1141
rect -2547 -1181 -2355 -1175
rect -2289 -1141 -2097 -1135
rect -2289 -1175 -2277 -1141
rect -2109 -1175 -2097 -1141
rect -2289 -1181 -2097 -1175
rect -2031 -1141 -1839 -1135
rect -2031 -1175 -2019 -1141
rect -1851 -1175 -1839 -1141
rect -2031 -1181 -1839 -1175
rect -1773 -1141 -1581 -1135
rect -1773 -1175 -1761 -1141
rect -1593 -1175 -1581 -1141
rect -1773 -1181 -1581 -1175
rect -1515 -1141 -1323 -1135
rect -1515 -1175 -1503 -1141
rect -1335 -1175 -1323 -1141
rect -1515 -1181 -1323 -1175
rect -1257 -1141 -1065 -1135
rect -1257 -1175 -1245 -1141
rect -1077 -1175 -1065 -1141
rect -1257 -1181 -1065 -1175
rect -999 -1141 -807 -1135
rect -999 -1175 -987 -1141
rect -819 -1175 -807 -1141
rect -999 -1181 -807 -1175
rect -741 -1141 -549 -1135
rect -741 -1175 -729 -1141
rect -561 -1175 -549 -1141
rect -741 -1181 -549 -1175
rect -483 -1141 -291 -1135
rect -483 -1175 -471 -1141
rect -303 -1175 -291 -1141
rect -483 -1181 -291 -1175
rect -225 -1141 -33 -1135
rect -225 -1175 -213 -1141
rect -45 -1175 -33 -1141
rect -225 -1181 -33 -1175
rect 33 -1141 225 -1135
rect 33 -1175 45 -1141
rect 213 -1175 225 -1141
rect 33 -1181 225 -1175
rect 291 -1141 483 -1135
rect 291 -1175 303 -1141
rect 471 -1175 483 -1141
rect 291 -1181 483 -1175
rect 549 -1141 741 -1135
rect 549 -1175 561 -1141
rect 729 -1175 741 -1141
rect 549 -1181 741 -1175
rect 807 -1141 999 -1135
rect 807 -1175 819 -1141
rect 987 -1175 999 -1141
rect 807 -1181 999 -1175
rect 1065 -1141 1257 -1135
rect 1065 -1175 1077 -1141
rect 1245 -1175 1257 -1141
rect 1065 -1181 1257 -1175
rect 1323 -1141 1515 -1135
rect 1323 -1175 1335 -1141
rect 1503 -1175 1515 -1141
rect 1323 -1181 1515 -1175
rect 1581 -1141 1773 -1135
rect 1581 -1175 1593 -1141
rect 1761 -1175 1773 -1141
rect 1581 -1181 1773 -1175
rect 1839 -1141 2031 -1135
rect 1839 -1175 1851 -1141
rect 2019 -1175 2031 -1141
rect 1839 -1181 2031 -1175
rect 2097 -1141 2289 -1135
rect 2097 -1175 2109 -1141
rect 2277 -1175 2289 -1141
rect 2097 -1181 2289 -1175
rect 2355 -1141 2547 -1135
rect 2355 -1175 2367 -1141
rect 2535 -1175 2547 -1141
rect 2355 -1181 2547 -1175
rect -2603 -1234 -2557 -1222
rect -2603 -1710 -2597 -1234
rect -2563 -1710 -2557 -1234
rect -2603 -1722 -2557 -1710
rect -2345 -1234 -2299 -1222
rect -2345 -1710 -2339 -1234
rect -2305 -1710 -2299 -1234
rect -2345 -1722 -2299 -1710
rect -2087 -1234 -2041 -1222
rect -2087 -1710 -2081 -1234
rect -2047 -1710 -2041 -1234
rect -2087 -1722 -2041 -1710
rect -1829 -1234 -1783 -1222
rect -1829 -1710 -1823 -1234
rect -1789 -1710 -1783 -1234
rect -1829 -1722 -1783 -1710
rect -1571 -1234 -1525 -1222
rect -1571 -1710 -1565 -1234
rect -1531 -1710 -1525 -1234
rect -1571 -1722 -1525 -1710
rect -1313 -1234 -1267 -1222
rect -1313 -1710 -1307 -1234
rect -1273 -1710 -1267 -1234
rect -1313 -1722 -1267 -1710
rect -1055 -1234 -1009 -1222
rect -1055 -1710 -1049 -1234
rect -1015 -1710 -1009 -1234
rect -1055 -1722 -1009 -1710
rect -797 -1234 -751 -1222
rect -797 -1710 -791 -1234
rect -757 -1710 -751 -1234
rect -797 -1722 -751 -1710
rect -539 -1234 -493 -1222
rect -539 -1710 -533 -1234
rect -499 -1710 -493 -1234
rect -539 -1722 -493 -1710
rect -281 -1234 -235 -1222
rect -281 -1710 -275 -1234
rect -241 -1710 -235 -1234
rect -281 -1722 -235 -1710
rect -23 -1234 23 -1222
rect -23 -1710 -17 -1234
rect 17 -1710 23 -1234
rect -23 -1722 23 -1710
rect 235 -1234 281 -1222
rect 235 -1710 241 -1234
rect 275 -1710 281 -1234
rect 235 -1722 281 -1710
rect 493 -1234 539 -1222
rect 493 -1710 499 -1234
rect 533 -1710 539 -1234
rect 493 -1722 539 -1710
rect 751 -1234 797 -1222
rect 751 -1710 757 -1234
rect 791 -1710 797 -1234
rect 751 -1722 797 -1710
rect 1009 -1234 1055 -1222
rect 1009 -1710 1015 -1234
rect 1049 -1710 1055 -1234
rect 1009 -1722 1055 -1710
rect 1267 -1234 1313 -1222
rect 1267 -1710 1273 -1234
rect 1307 -1710 1313 -1234
rect 1267 -1722 1313 -1710
rect 1525 -1234 1571 -1222
rect 1525 -1710 1531 -1234
rect 1565 -1710 1571 -1234
rect 1525 -1722 1571 -1710
rect 1783 -1234 1829 -1222
rect 1783 -1710 1789 -1234
rect 1823 -1710 1829 -1234
rect 1783 -1722 1829 -1710
rect 2041 -1234 2087 -1222
rect 2041 -1710 2047 -1234
rect 2081 -1710 2087 -1234
rect 2041 -1722 2087 -1710
rect 2299 -1234 2345 -1222
rect 2299 -1710 2305 -1234
rect 2339 -1710 2345 -1234
rect 2299 -1722 2345 -1710
rect 2557 -1234 2603 -1222
rect 2557 -1710 2563 -1234
rect 2597 -1710 2603 -1234
rect 2557 -1722 2603 -1710
rect -2547 -1769 -2355 -1763
rect -2547 -1803 -2535 -1769
rect -2367 -1803 -2355 -1769
rect -2547 -1809 -2355 -1803
rect -2289 -1769 -2097 -1763
rect -2289 -1803 -2277 -1769
rect -2109 -1803 -2097 -1769
rect -2289 -1809 -2097 -1803
rect -2031 -1769 -1839 -1763
rect -2031 -1803 -2019 -1769
rect -1851 -1803 -1839 -1769
rect -2031 -1809 -1839 -1803
rect -1773 -1769 -1581 -1763
rect -1773 -1803 -1761 -1769
rect -1593 -1803 -1581 -1769
rect -1773 -1809 -1581 -1803
rect -1515 -1769 -1323 -1763
rect -1515 -1803 -1503 -1769
rect -1335 -1803 -1323 -1769
rect -1515 -1809 -1323 -1803
rect -1257 -1769 -1065 -1763
rect -1257 -1803 -1245 -1769
rect -1077 -1803 -1065 -1769
rect -1257 -1809 -1065 -1803
rect -999 -1769 -807 -1763
rect -999 -1803 -987 -1769
rect -819 -1803 -807 -1769
rect -999 -1809 -807 -1803
rect -741 -1769 -549 -1763
rect -741 -1803 -729 -1769
rect -561 -1803 -549 -1769
rect -741 -1809 -549 -1803
rect -483 -1769 -291 -1763
rect -483 -1803 -471 -1769
rect -303 -1803 -291 -1769
rect -483 -1809 -291 -1803
rect -225 -1769 -33 -1763
rect -225 -1803 -213 -1769
rect -45 -1803 -33 -1769
rect -225 -1809 -33 -1803
rect 33 -1769 225 -1763
rect 33 -1803 45 -1769
rect 213 -1803 225 -1769
rect 33 -1809 225 -1803
rect 291 -1769 483 -1763
rect 291 -1803 303 -1769
rect 471 -1803 483 -1769
rect 291 -1809 483 -1803
rect 549 -1769 741 -1763
rect 549 -1803 561 -1769
rect 729 -1803 741 -1769
rect 549 -1809 741 -1803
rect 807 -1769 999 -1763
rect 807 -1803 819 -1769
rect 987 -1803 999 -1769
rect 807 -1809 999 -1803
rect 1065 -1769 1257 -1763
rect 1065 -1803 1077 -1769
rect 1245 -1803 1257 -1769
rect 1065 -1809 1257 -1803
rect 1323 -1769 1515 -1763
rect 1323 -1803 1335 -1769
rect 1503 -1803 1515 -1769
rect 1323 -1809 1515 -1803
rect 1581 -1769 1773 -1763
rect 1581 -1803 1593 -1769
rect 1761 -1803 1773 -1769
rect 1581 -1809 1773 -1803
rect 1839 -1769 2031 -1763
rect 1839 -1803 1851 -1769
rect 2019 -1803 2031 -1769
rect 1839 -1809 2031 -1803
rect 2097 -1769 2289 -1763
rect 2097 -1803 2109 -1769
rect 2277 -1803 2289 -1769
rect 2097 -1809 2289 -1803
rect 2355 -1769 2547 -1763
rect 2355 -1803 2367 -1769
rect 2535 -1803 2547 -1769
rect 2355 -1809 2547 -1803
rect -2547 -1877 -2355 -1871
rect -2547 -1911 -2535 -1877
rect -2367 -1911 -2355 -1877
rect -2547 -1917 -2355 -1911
rect -2289 -1877 -2097 -1871
rect -2289 -1911 -2277 -1877
rect -2109 -1911 -2097 -1877
rect -2289 -1917 -2097 -1911
rect -2031 -1877 -1839 -1871
rect -2031 -1911 -2019 -1877
rect -1851 -1911 -1839 -1877
rect -2031 -1917 -1839 -1911
rect -1773 -1877 -1581 -1871
rect -1773 -1911 -1761 -1877
rect -1593 -1911 -1581 -1877
rect -1773 -1917 -1581 -1911
rect -1515 -1877 -1323 -1871
rect -1515 -1911 -1503 -1877
rect -1335 -1911 -1323 -1877
rect -1515 -1917 -1323 -1911
rect -1257 -1877 -1065 -1871
rect -1257 -1911 -1245 -1877
rect -1077 -1911 -1065 -1877
rect -1257 -1917 -1065 -1911
rect -999 -1877 -807 -1871
rect -999 -1911 -987 -1877
rect -819 -1911 -807 -1877
rect -999 -1917 -807 -1911
rect -741 -1877 -549 -1871
rect -741 -1911 -729 -1877
rect -561 -1911 -549 -1877
rect -741 -1917 -549 -1911
rect -483 -1877 -291 -1871
rect -483 -1911 -471 -1877
rect -303 -1911 -291 -1877
rect -483 -1917 -291 -1911
rect -225 -1877 -33 -1871
rect -225 -1911 -213 -1877
rect -45 -1911 -33 -1877
rect -225 -1917 -33 -1911
rect 33 -1877 225 -1871
rect 33 -1911 45 -1877
rect 213 -1911 225 -1877
rect 33 -1917 225 -1911
rect 291 -1877 483 -1871
rect 291 -1911 303 -1877
rect 471 -1911 483 -1877
rect 291 -1917 483 -1911
rect 549 -1877 741 -1871
rect 549 -1911 561 -1877
rect 729 -1911 741 -1877
rect 549 -1917 741 -1911
rect 807 -1877 999 -1871
rect 807 -1911 819 -1877
rect 987 -1911 999 -1877
rect 807 -1917 999 -1911
rect 1065 -1877 1257 -1871
rect 1065 -1911 1077 -1877
rect 1245 -1911 1257 -1877
rect 1065 -1917 1257 -1911
rect 1323 -1877 1515 -1871
rect 1323 -1911 1335 -1877
rect 1503 -1911 1515 -1877
rect 1323 -1917 1515 -1911
rect 1581 -1877 1773 -1871
rect 1581 -1911 1593 -1877
rect 1761 -1911 1773 -1877
rect 1581 -1917 1773 -1911
rect 1839 -1877 2031 -1871
rect 1839 -1911 1851 -1877
rect 2019 -1911 2031 -1877
rect 1839 -1917 2031 -1911
rect 2097 -1877 2289 -1871
rect 2097 -1911 2109 -1877
rect 2277 -1911 2289 -1877
rect 2097 -1917 2289 -1911
rect 2355 -1877 2547 -1871
rect 2355 -1911 2367 -1877
rect 2535 -1911 2547 -1877
rect 2355 -1917 2547 -1911
rect -2603 -1970 -2557 -1958
rect -2603 -2446 -2597 -1970
rect -2563 -2446 -2557 -1970
rect -2603 -2458 -2557 -2446
rect -2345 -1970 -2299 -1958
rect -2345 -2446 -2339 -1970
rect -2305 -2446 -2299 -1970
rect -2345 -2458 -2299 -2446
rect -2087 -1970 -2041 -1958
rect -2087 -2446 -2081 -1970
rect -2047 -2446 -2041 -1970
rect -2087 -2458 -2041 -2446
rect -1829 -1970 -1783 -1958
rect -1829 -2446 -1823 -1970
rect -1789 -2446 -1783 -1970
rect -1829 -2458 -1783 -2446
rect -1571 -1970 -1525 -1958
rect -1571 -2446 -1565 -1970
rect -1531 -2446 -1525 -1970
rect -1571 -2458 -1525 -2446
rect -1313 -1970 -1267 -1958
rect -1313 -2446 -1307 -1970
rect -1273 -2446 -1267 -1970
rect -1313 -2458 -1267 -2446
rect -1055 -1970 -1009 -1958
rect -1055 -2446 -1049 -1970
rect -1015 -2446 -1009 -1970
rect -1055 -2458 -1009 -2446
rect -797 -1970 -751 -1958
rect -797 -2446 -791 -1970
rect -757 -2446 -751 -1970
rect -797 -2458 -751 -2446
rect -539 -1970 -493 -1958
rect -539 -2446 -533 -1970
rect -499 -2446 -493 -1970
rect -539 -2458 -493 -2446
rect -281 -1970 -235 -1958
rect -281 -2446 -275 -1970
rect -241 -2446 -235 -1970
rect -281 -2458 -235 -2446
rect -23 -1970 23 -1958
rect -23 -2446 -17 -1970
rect 17 -2446 23 -1970
rect -23 -2458 23 -2446
rect 235 -1970 281 -1958
rect 235 -2446 241 -1970
rect 275 -2446 281 -1970
rect 235 -2458 281 -2446
rect 493 -1970 539 -1958
rect 493 -2446 499 -1970
rect 533 -2446 539 -1970
rect 493 -2458 539 -2446
rect 751 -1970 797 -1958
rect 751 -2446 757 -1970
rect 791 -2446 797 -1970
rect 751 -2458 797 -2446
rect 1009 -1970 1055 -1958
rect 1009 -2446 1015 -1970
rect 1049 -2446 1055 -1970
rect 1009 -2458 1055 -2446
rect 1267 -1970 1313 -1958
rect 1267 -2446 1273 -1970
rect 1307 -2446 1313 -1970
rect 1267 -2458 1313 -2446
rect 1525 -1970 1571 -1958
rect 1525 -2446 1531 -1970
rect 1565 -2446 1571 -1970
rect 1525 -2458 1571 -2446
rect 1783 -1970 1829 -1958
rect 1783 -2446 1789 -1970
rect 1823 -2446 1829 -1970
rect 1783 -2458 1829 -2446
rect 2041 -1970 2087 -1958
rect 2041 -2446 2047 -1970
rect 2081 -2446 2087 -1970
rect 2041 -2458 2087 -2446
rect 2299 -1970 2345 -1958
rect 2299 -2446 2305 -1970
rect 2339 -2446 2345 -1970
rect 2299 -2458 2345 -2446
rect 2557 -1970 2603 -1958
rect 2557 -2446 2563 -1970
rect 2597 -2446 2603 -1970
rect 2557 -2458 2603 -2446
rect -2547 -2505 -2355 -2499
rect -2547 -2539 -2535 -2505
rect -2367 -2539 -2355 -2505
rect -2547 -2545 -2355 -2539
rect -2289 -2505 -2097 -2499
rect -2289 -2539 -2277 -2505
rect -2109 -2539 -2097 -2505
rect -2289 -2545 -2097 -2539
rect -2031 -2505 -1839 -2499
rect -2031 -2539 -2019 -2505
rect -1851 -2539 -1839 -2505
rect -2031 -2545 -1839 -2539
rect -1773 -2505 -1581 -2499
rect -1773 -2539 -1761 -2505
rect -1593 -2539 -1581 -2505
rect -1773 -2545 -1581 -2539
rect -1515 -2505 -1323 -2499
rect -1515 -2539 -1503 -2505
rect -1335 -2539 -1323 -2505
rect -1515 -2545 -1323 -2539
rect -1257 -2505 -1065 -2499
rect -1257 -2539 -1245 -2505
rect -1077 -2539 -1065 -2505
rect -1257 -2545 -1065 -2539
rect -999 -2505 -807 -2499
rect -999 -2539 -987 -2505
rect -819 -2539 -807 -2505
rect -999 -2545 -807 -2539
rect -741 -2505 -549 -2499
rect -741 -2539 -729 -2505
rect -561 -2539 -549 -2505
rect -741 -2545 -549 -2539
rect -483 -2505 -291 -2499
rect -483 -2539 -471 -2505
rect -303 -2539 -291 -2505
rect -483 -2545 -291 -2539
rect -225 -2505 -33 -2499
rect -225 -2539 -213 -2505
rect -45 -2539 -33 -2505
rect -225 -2545 -33 -2539
rect 33 -2505 225 -2499
rect 33 -2539 45 -2505
rect 213 -2539 225 -2505
rect 33 -2545 225 -2539
rect 291 -2505 483 -2499
rect 291 -2539 303 -2505
rect 471 -2539 483 -2505
rect 291 -2545 483 -2539
rect 549 -2505 741 -2499
rect 549 -2539 561 -2505
rect 729 -2539 741 -2505
rect 549 -2545 741 -2539
rect 807 -2505 999 -2499
rect 807 -2539 819 -2505
rect 987 -2539 999 -2505
rect 807 -2545 999 -2539
rect 1065 -2505 1257 -2499
rect 1065 -2539 1077 -2505
rect 1245 -2539 1257 -2505
rect 1065 -2545 1257 -2539
rect 1323 -2505 1515 -2499
rect 1323 -2539 1335 -2505
rect 1503 -2539 1515 -2505
rect 1323 -2545 1515 -2539
rect 1581 -2505 1773 -2499
rect 1581 -2539 1593 -2505
rect 1761 -2539 1773 -2505
rect 1581 -2545 1773 -2539
rect 1839 -2505 2031 -2499
rect 1839 -2539 1851 -2505
rect 2019 -2539 2031 -2505
rect 1839 -2545 2031 -2539
rect 2097 -2505 2289 -2499
rect 2097 -2539 2109 -2505
rect 2277 -2539 2289 -2505
rect 2097 -2545 2289 -2539
rect 2355 -2505 2547 -2499
rect 2355 -2539 2367 -2505
rect 2535 -2539 2547 -2505
rect 2355 -2545 2547 -2539
<< properties >>
string FIXED_BBOX -2694 -2624 2694 2624
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.5 l 1.0 m 7 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
