magic
tech sky130A
magscale 1 2
timestamp 1713391016
<< error_s >>
rect 20758 7946 20816 7952
rect 20950 7946 21008 7952
rect 21142 7946 21200 7952
rect 21334 7946 21392 7952
rect 21526 7946 21584 7952
rect 20758 7912 20770 7946
rect 20950 7912 20962 7946
rect 21142 7912 21154 7946
rect 21334 7912 21346 7946
rect 21526 7912 21538 7946
rect 20758 7906 20816 7912
rect 20950 7906 21008 7912
rect 21142 7906 21200 7912
rect 21334 7906 21392 7912
rect 21526 7906 21584 7912
rect 20662 6818 20720 6824
rect 20854 6818 20912 6824
rect 21046 6818 21104 6824
rect 21238 6818 21296 6824
rect 21430 6818 21488 6824
rect 20662 6784 20674 6818
rect 20854 6784 20866 6818
rect 21046 6784 21058 6818
rect 21238 6784 21250 6818
rect 21430 6784 21442 6818
rect 20662 6778 20720 6784
rect 20854 6778 20912 6784
rect 21046 6778 21104 6784
rect 21238 6778 21296 6784
rect 21430 6778 21488 6784
rect 20650 6178 20708 6184
rect 20842 6178 20900 6184
rect 21034 6178 21092 6184
rect 21226 6178 21284 6184
rect 21418 6178 21476 6184
rect 20650 6144 20662 6178
rect 20842 6144 20854 6178
rect 21034 6144 21046 6178
rect 21226 6144 21238 6178
rect 21418 6144 21430 6178
rect 20650 6138 20708 6144
rect 20842 6138 20900 6144
rect 21034 6138 21092 6144
rect 21226 6138 21284 6144
rect 21418 6138 21476 6144
rect 20746 5268 20804 5274
rect 20938 5268 20996 5274
rect 21130 5268 21188 5274
rect 21322 5268 21380 5274
rect 21514 5268 21572 5274
rect 20746 5234 20758 5268
rect 20938 5234 20950 5268
rect 21130 5234 21142 5268
rect 21322 5234 21334 5268
rect 21514 5234 21526 5268
rect 20746 5228 20804 5234
rect 20938 5228 20996 5234
rect 21130 5228 21188 5234
rect 21322 5228 21380 5234
rect 21514 5228 21572 5234
rect 20746 5160 20804 5166
rect 20938 5160 20996 5166
rect 21130 5160 21188 5166
rect 21322 5160 21380 5166
rect 21514 5160 21572 5166
rect 20746 5126 20758 5160
rect 20938 5126 20950 5160
rect 21130 5126 21142 5160
rect 21322 5126 21334 5160
rect 21514 5126 21526 5160
rect 20746 5120 20804 5126
rect 20938 5120 20996 5126
rect 21130 5120 21188 5126
rect 21322 5120 21380 5126
rect 21514 5120 21572 5126
rect 20650 4250 20708 4256
rect 20842 4250 20900 4256
rect 21034 4250 21092 4256
rect 21226 4250 21284 4256
rect 21418 4250 21476 4256
rect 20650 4216 20662 4250
rect 20842 4216 20854 4250
rect 21034 4216 21046 4250
rect 21226 4216 21238 4250
rect 21418 4216 21430 4250
rect 20650 4210 20708 4216
rect 20842 4210 20900 4216
rect 21034 4210 21092 4216
rect 21226 4210 21284 4216
rect 21418 4210 21476 4216
<< pwell >>
rect 1872 7070 1982 7542
rect 2684 7472 2800 7944
rect 5588 7716 7106 7774
rect 5272 7484 5532 7544
rect 5588 7398 7106 7456
rect 5588 7300 7106 7358
rect 5274 7066 5532 7128
rect 5588 6982 7106 7040
rect 5588 6884 7106 6942
rect 5274 6654 5528 6708
rect 5588 6566 7106 6624
rect 5588 6462 7106 6520
rect 5588 6146 7106 6204
rect 5594 6046 7112 6104
rect 5588 5730 7106 5788
rect 2564 2372 2632 2528
rect 3484 2372 3552 2528
rect 4398 2372 4466 2528
rect 5314 2372 5382 2528
<< viali >>
rect 4352 9918 4562 9988
rect 6330 9916 6522 9984
rect 8164 9936 8432 10006
rect 12314 9934 12618 10008
rect 14222 9936 14510 10006
rect 18376 9932 18668 10008
rect 20274 9878 20448 9954
rect 21366 9880 21528 9956
rect 4556 5626 4794 5684
rect 6034 5624 6276 5686
rect 1078 4942 1242 4998
rect 1472 4942 1636 4998
rect 1866 4942 2030 4998
rect 2258 4942 2428 5000
rect 2670 4942 2834 5000
rect 3062 4942 3224 5000
rect 1068 3292 1142 3556
rect 8684 3202 9426 3266
rect 2038 2042 2246 2134
rect 4814 2046 5046 2134
rect 7516 2052 7754 2138
rect 10260 2052 10500 2136
rect 12758 2052 12986 2138
rect 15548 2054 15776 2136
rect 17912 2060 18164 2136
rect 20726 2056 20964 2136
<< metal1 >>
rect 30 10348 22606 10794
rect 546 10136 752 10348
rect 3508 10178 3600 10348
rect 3502 10086 3508 10178
rect 3600 10086 3606 10178
rect 546 9924 752 9930
rect 4312 9988 4604 10348
rect 4312 9918 4352 9988
rect 4562 9918 4604 9988
rect 4312 9908 4604 9918
rect 6276 9984 6568 10348
rect 7264 10179 7359 10348
rect 7258 10084 7264 10179
rect 7359 10084 7365 10179
rect 6276 9916 6330 9984
rect 6522 9916 6568 9984
rect 8088 10006 8492 10348
rect 8088 9936 8164 10006
rect 8432 9936 8492 10006
rect 8088 9922 8492 9936
rect 12264 10008 12668 10348
rect 13417 10171 13552 10348
rect 13411 10036 13417 10171
rect 13552 10036 13558 10171
rect 12264 9934 12314 10008
rect 12618 9934 12668 10008
rect 12264 9920 12668 9934
rect 14158 10006 14562 10348
rect 14158 9936 14222 10006
rect 14510 9936 14562 10006
rect 14158 9924 14562 9936
rect 18324 10008 18728 10348
rect 18324 9932 18376 10008
rect 18668 9932 18728 10008
rect 18324 9922 18728 9932
rect 20240 9954 20478 10348
rect 6276 9906 6568 9916
rect 3830 9816 7048 9876
rect 7898 9840 19096 9890
rect 20240 9878 20274 9954
rect 20448 9878 20478 9954
rect 20240 9870 20478 9878
rect 21332 9956 21570 10348
rect 21332 9880 21366 9956
rect 21528 9880 21570 9956
rect 21332 9866 21570 9880
rect 3768 9718 3778 9774
rect 3840 9718 3850 9774
rect 4282 9720 4292 9776
rect 4354 9720 4364 9776
rect 4800 9722 4810 9778
rect 4872 9722 4882 9778
rect 4024 9592 4034 9652
rect 4098 9592 4108 9652
rect 4540 9592 4550 9652
rect 4614 9592 4624 9652
rect 5056 9592 5066 9652
rect 5130 9592 5140 9652
rect 5275 9640 5329 9646
rect 5370 9640 5476 9816
rect 5980 9722 5990 9778
rect 6052 9722 6062 9778
rect 6498 9722 6508 9778
rect 6570 9722 6580 9778
rect 7014 9722 7024 9778
rect 7086 9722 7096 9778
rect 7834 9712 7844 9798
rect 7912 9712 7922 9798
rect 8352 9712 8362 9798
rect 8430 9712 8440 9798
rect 8868 9712 8878 9798
rect 8946 9712 8956 9798
rect 9384 9712 9394 9798
rect 9462 9712 9472 9798
rect 9900 9712 9910 9798
rect 9978 9712 9988 9798
rect 10416 9712 10426 9798
rect 10494 9712 10504 9798
rect 10932 9712 10942 9798
rect 11010 9712 11020 9798
rect 11448 9712 11458 9798
rect 11526 9712 11536 9798
rect 11962 9712 11972 9798
rect 12040 9712 12050 9798
rect 12480 9712 12490 9798
rect 12558 9712 12568 9798
rect 12996 9712 13006 9798
rect 13074 9712 13084 9798
rect 5329 9586 5476 9640
rect 5275 9580 5329 9586
rect 5370 9548 5476 9586
rect 5724 9584 5734 9644
rect 5798 9584 5808 9644
rect 6238 9584 6248 9644
rect 6312 9584 6322 9644
rect 6756 9584 6766 9644
rect 6830 9584 6840 9644
rect 3830 9488 7048 9548
rect 13376 9262 13592 9840
rect 13908 9712 13918 9798
rect 13986 9712 13996 9798
rect 14422 9712 14432 9798
rect 14500 9712 14510 9798
rect 14938 9712 14948 9798
rect 15016 9712 15026 9798
rect 15454 9712 15464 9798
rect 15532 9712 15542 9798
rect 15972 9712 15982 9798
rect 16050 9712 16060 9798
rect 16486 9712 16496 9798
rect 16564 9712 16574 9798
rect 17004 9712 17014 9798
rect 17082 9712 17092 9798
rect 17518 9712 17528 9798
rect 17596 9712 17606 9798
rect 18036 9712 18046 9798
rect 18114 9712 18124 9798
rect 18550 9712 18560 9798
rect 18628 9712 18638 9798
rect 19068 9712 19078 9798
rect 19146 9712 19156 9798
rect 7900 9212 19098 9262
rect 13376 9152 13592 9212
rect 7900 9102 19098 9152
rect 7834 8974 7844 9060
rect 7912 8974 7922 9060
rect 8350 8974 8360 9060
rect 8428 8974 8438 9060
rect 8868 8974 8878 9060
rect 8946 8974 8956 9060
rect 9382 8974 9392 9060
rect 9460 8974 9470 9060
rect 9898 8974 9908 9060
rect 9976 8974 9986 9060
rect 10414 8974 10424 9060
rect 10492 8974 10502 9060
rect 10930 8974 10940 9060
rect 11008 8974 11018 9060
rect 11446 8976 11456 9062
rect 11524 8976 11534 9062
rect 11962 8976 11972 9062
rect 12040 8976 12050 9062
rect 12478 8976 12488 9062
rect 12556 8976 12566 9062
rect 12996 8976 13006 9062
rect 13074 8976 13084 9062
rect 13376 8528 13592 9102
rect 13908 8976 13918 9062
rect 13986 8976 13996 9062
rect 14422 8976 14432 9062
rect 14500 8976 14510 9062
rect 14938 8976 14948 9062
rect 15016 8976 15026 9062
rect 15456 8976 15466 9062
rect 15534 8976 15544 9062
rect 15968 8976 15978 9062
rect 16046 8976 16056 9062
rect 16486 8972 16496 9058
rect 16564 8972 16574 9058
rect 17002 8972 17012 9058
rect 17080 8972 17090 9058
rect 17516 8972 17526 9058
rect 17594 8972 17604 9058
rect 18034 8972 18044 9058
rect 18112 8972 18122 9058
rect 18552 8972 18562 9058
rect 18630 8972 18640 9058
rect 19068 8972 19078 9058
rect 19146 8972 19156 9058
rect 102 8284 3830 8484
rect 7900 8478 19098 8528
rect 13376 8418 13592 8478
rect 7900 8368 19098 8418
rect 3630 8096 3830 8284
rect 7834 8246 7844 8332
rect 7912 8246 7922 8332
rect 8350 8246 8360 8332
rect 8428 8246 8438 8332
rect 8866 8246 8876 8332
rect 8944 8246 8954 8332
rect 9382 8246 9392 8332
rect 9460 8246 9470 8332
rect 9898 8246 9908 8332
rect 9976 8246 9986 8332
rect 10414 8246 10424 8332
rect 10492 8246 10502 8332
rect 10930 8246 10940 8332
rect 11008 8246 11018 8332
rect 11446 8246 11456 8332
rect 11524 8246 11534 8332
rect 11962 8246 11972 8332
rect 12040 8246 12050 8332
rect 12478 8246 12488 8332
rect 12556 8246 12566 8332
rect 12994 8246 13004 8332
rect 13072 8246 13082 8332
rect 2293 7542 2403 7941
rect 1128 7436 1610 7536
rect 540 6937 546 7143
rect 752 6937 758 7143
rect 1128 7074 1222 7436
rect 1510 7080 1610 7436
rect 1872 7432 2403 7542
rect 2684 7828 3202 7944
rect 2684 7472 2800 7828
rect 3086 7450 3202 7828
rect 3658 7774 3803 8096
rect 13376 7792 13592 8368
rect 13908 8244 13918 8330
rect 13986 8244 13996 8330
rect 14420 8244 14430 8330
rect 14498 8244 14508 8330
rect 14938 8244 14948 8330
rect 15016 8244 15026 8330
rect 15454 8244 15464 8330
rect 15532 8244 15542 8330
rect 15970 8244 15980 8330
rect 16048 8244 16058 8330
rect 16486 8244 16496 8330
rect 16564 8244 16574 8330
rect 17002 8244 17012 8330
rect 17080 8244 17090 8330
rect 17518 8244 17528 8330
rect 17596 8244 17606 8330
rect 18034 8244 18044 8330
rect 18112 8244 18122 8330
rect 18550 8244 18560 8330
rect 18628 8244 18638 8330
rect 19066 8244 19076 8330
rect 19144 8244 19154 8330
rect 3658 7716 5226 7774
rect 5588 7716 7106 7774
rect 7900 7742 19098 7792
rect 3658 7714 3803 7716
rect 3708 7456 3766 7714
rect 4020 7626 4030 7686
rect 4094 7626 4104 7686
rect 4254 7626 4264 7686
rect 4328 7626 4338 7686
rect 4490 7626 4500 7686
rect 4564 7626 4574 7686
rect 4726 7626 4736 7686
rect 4800 7626 4810 7686
rect 4962 7626 4972 7686
rect 5036 7626 5046 7686
rect 5198 7626 5208 7686
rect 5272 7626 5282 7686
rect 5526 7626 5536 7684
rect 5600 7626 5610 7684
rect 5762 7626 5772 7684
rect 5836 7626 5846 7684
rect 5998 7626 6008 7684
rect 6072 7626 6082 7684
rect 6234 7626 6244 7684
rect 6308 7626 6318 7684
rect 6470 7626 6480 7684
rect 6544 7626 6554 7684
rect 6706 7626 6716 7684
rect 6780 7626 6790 7684
rect 4134 7490 4144 7550
rect 4214 7490 4224 7550
rect 4370 7492 4380 7552
rect 4450 7492 4460 7552
rect 4606 7492 4616 7552
rect 4686 7492 4696 7552
rect 4840 7492 4850 7552
rect 4920 7492 4930 7552
rect 5078 7492 5088 7552
rect 5158 7492 5168 7552
rect 5646 7492 5656 7552
rect 5716 7492 5726 7552
rect 5882 7492 5892 7552
rect 5952 7492 5962 7552
rect 6118 7492 6128 7552
rect 6188 7492 6198 7552
rect 6354 7492 6364 7552
rect 6424 7492 6434 7552
rect 6590 7492 6600 7552
rect 6660 7492 6670 7552
rect 7045 7456 7103 7716
rect 13376 7682 13592 7742
rect 7900 7632 19098 7682
rect 7834 7504 7844 7590
rect 7912 7504 7922 7590
rect 8350 7504 8360 7590
rect 8428 7504 8438 7590
rect 8866 7504 8876 7590
rect 8944 7504 8954 7590
rect 9382 7504 9392 7590
rect 9460 7504 9470 7590
rect 9898 7504 9908 7590
rect 9976 7504 9986 7590
rect 10414 7504 10424 7590
rect 10492 7504 10502 7590
rect 10930 7504 10940 7590
rect 11008 7504 11018 7590
rect 11446 7504 11456 7590
rect 11524 7504 11534 7590
rect 11964 7504 11974 7590
rect 12042 7504 12052 7590
rect 12480 7504 12490 7590
rect 12558 7504 12568 7590
rect 12996 7504 13006 7590
rect 13074 7504 13084 7590
rect 1872 7070 1982 7432
rect 3708 7398 5226 7456
rect 5588 7398 7106 7456
rect 3708 7358 3766 7398
rect 7045 7358 7103 7398
rect 3708 7300 5226 7358
rect 5588 7300 7106 7358
rect 3708 7040 3766 7300
rect 4018 7208 4028 7268
rect 4092 7208 4102 7268
rect 4254 7208 4264 7268
rect 4328 7208 4338 7268
rect 4490 7208 4500 7268
rect 4564 7208 4574 7268
rect 4726 7208 4736 7268
rect 4800 7208 4810 7268
rect 4962 7208 4972 7268
rect 5036 7208 5046 7268
rect 5200 7208 5210 7268
rect 5274 7208 5284 7268
rect 5526 7208 5536 7266
rect 5600 7208 5610 7266
rect 5762 7208 5772 7266
rect 5836 7208 5846 7266
rect 5998 7208 6008 7266
rect 6072 7208 6082 7266
rect 6234 7208 6244 7266
rect 6308 7208 6318 7266
rect 6470 7208 6480 7266
rect 6544 7208 6554 7266
rect 6706 7208 6716 7266
rect 6780 7208 6790 7266
rect 4132 7076 4142 7136
rect 4212 7076 4222 7136
rect 4370 7076 4380 7136
rect 4450 7076 4460 7136
rect 4606 7076 4616 7136
rect 4686 7076 4696 7136
rect 4842 7076 4852 7136
rect 4922 7076 4932 7136
rect 5078 7076 5088 7136
rect 5158 7076 5168 7136
rect 5646 7072 5656 7132
rect 5716 7072 5726 7132
rect 5882 7072 5892 7132
rect 5952 7072 5962 7132
rect 6118 7072 6128 7132
rect 6188 7072 6198 7132
rect 6354 7072 6364 7132
rect 6424 7072 6434 7132
rect 6590 7072 6600 7132
rect 6660 7072 6670 7132
rect 7045 7040 7103 7300
rect 13376 7056 13592 7632
rect 13906 7504 13916 7590
rect 13984 7504 13994 7590
rect 14422 7504 14432 7590
rect 14500 7504 14510 7590
rect 14938 7504 14948 7590
rect 15016 7504 15026 7590
rect 15454 7504 15464 7590
rect 15532 7504 15542 7590
rect 15970 7504 15980 7590
rect 16048 7504 16058 7590
rect 16486 7504 16496 7590
rect 16564 7504 16574 7590
rect 17002 7504 17012 7590
rect 17080 7504 17090 7590
rect 17518 7504 17528 7590
rect 17596 7504 17606 7590
rect 18034 7504 18044 7590
rect 18112 7504 18122 7590
rect 18550 7504 18560 7590
rect 18628 7504 18638 7590
rect 19068 7504 19078 7590
rect 19146 7504 19156 7590
rect 3708 6982 5226 7040
rect 5588 6982 7106 7040
rect 7900 7006 19098 7056
rect 3708 6942 3766 6982
rect 7045 6942 7103 6982
rect 13376 6946 13592 7006
rect 546 5338 752 6937
rect 3708 6884 5226 6942
rect 5588 6884 7106 6942
rect 7900 6896 19098 6946
rect 3708 6624 3766 6884
rect 4018 6788 4028 6848
rect 4092 6788 4102 6848
rect 4254 6790 4264 6850
rect 4328 6790 4338 6850
rect 4492 6790 4502 6850
rect 4566 6790 4576 6850
rect 4726 6790 4736 6850
rect 4800 6790 4810 6850
rect 4962 6790 4972 6850
rect 5036 6790 5046 6850
rect 5198 6790 5208 6850
rect 5272 6790 5282 6850
rect 5526 6792 5536 6850
rect 5600 6792 5610 6850
rect 5762 6792 5772 6850
rect 5836 6792 5846 6850
rect 6000 6792 6010 6850
rect 6074 6792 6084 6850
rect 6234 6792 6244 6850
rect 6308 6792 6318 6850
rect 6470 6792 6480 6850
rect 6544 6792 6554 6850
rect 6706 6794 6716 6852
rect 6780 6794 6790 6852
rect 4132 6656 4142 6716
rect 4212 6656 4222 6716
rect 4370 6656 4380 6716
rect 4450 6656 4460 6716
rect 4606 6656 4616 6716
rect 4686 6656 4696 6716
rect 4842 6656 4852 6716
rect 4922 6656 4932 6716
rect 5080 6656 5090 6716
rect 5160 6656 5170 6716
rect 5646 6660 5656 6720
rect 5716 6660 5726 6720
rect 5882 6660 5892 6720
rect 5952 6660 5962 6720
rect 6118 6660 6128 6720
rect 6188 6660 6198 6720
rect 6354 6660 6364 6720
rect 6424 6660 6434 6720
rect 6590 6660 6600 6720
rect 6660 6660 6670 6720
rect 7045 6624 7103 6884
rect 7834 6776 7844 6862
rect 7912 6776 7922 6862
rect 8350 6776 8360 6862
rect 8428 6776 8438 6862
rect 8864 6776 8874 6862
rect 8942 6776 8952 6862
rect 9382 6776 9392 6862
rect 9460 6776 9470 6862
rect 9898 6776 9908 6862
rect 9976 6776 9986 6862
rect 10414 6776 10424 6862
rect 10492 6776 10502 6862
rect 10930 6776 10940 6862
rect 11008 6776 11018 6862
rect 11446 6776 11456 6862
rect 11524 6776 11534 6862
rect 11962 6776 11972 6862
rect 12040 6776 12050 6862
rect 12478 6776 12488 6862
rect 12556 6776 12566 6862
rect 12996 6776 13006 6862
rect 13074 6776 13084 6862
rect 3708 6566 5226 6624
rect 5588 6566 7106 6624
rect 3708 6520 3766 6566
rect 7045 6520 7103 6566
rect 3708 6462 5226 6520
rect 5588 6462 7106 6520
rect 3708 6204 3766 6462
rect 4018 6374 4028 6434
rect 4092 6374 4102 6434
rect 4254 6374 4264 6434
rect 4328 6374 4338 6434
rect 4490 6374 4500 6434
rect 4564 6374 4574 6434
rect 4726 6374 4736 6434
rect 4800 6374 4810 6434
rect 4962 6374 4972 6434
rect 5036 6374 5046 6434
rect 5198 6374 5208 6434
rect 5272 6374 5282 6434
rect 5526 6376 5536 6434
rect 5600 6376 5610 6434
rect 5762 6376 5772 6434
rect 5836 6376 5846 6434
rect 5998 6376 6008 6434
rect 6072 6376 6082 6434
rect 6234 6376 6244 6434
rect 6308 6376 6318 6434
rect 6470 6376 6480 6434
rect 6544 6376 6554 6434
rect 6706 6376 6716 6434
rect 6780 6376 6790 6434
rect 4134 6240 4144 6300
rect 4214 6240 4224 6300
rect 4370 6240 4380 6300
rect 4450 6240 4460 6300
rect 4606 6240 4616 6300
rect 4686 6240 4696 6300
rect 4842 6240 4852 6300
rect 4922 6240 4932 6300
rect 5078 6240 5088 6300
rect 5158 6240 5168 6300
rect 5646 6244 5656 6304
rect 5716 6244 5726 6304
rect 5882 6244 5892 6304
rect 5952 6244 5962 6304
rect 6118 6244 6128 6304
rect 6188 6244 6198 6304
rect 6354 6244 6364 6304
rect 6424 6244 6434 6304
rect 6590 6244 6600 6304
rect 6660 6244 6670 6304
rect 7045 6204 7103 6462
rect 13376 6320 13592 6896
rect 13906 6776 13916 6862
rect 13984 6776 13994 6862
rect 14420 6776 14430 6862
rect 14498 6776 14508 6862
rect 14938 6776 14948 6862
rect 15016 6776 15026 6862
rect 15454 6776 15464 6862
rect 15532 6776 15542 6862
rect 15970 6776 15980 6862
rect 16048 6776 16058 6862
rect 16488 6776 16498 6862
rect 16566 6776 16576 6862
rect 17000 6776 17010 6862
rect 17078 6776 17088 6862
rect 17518 6776 17528 6862
rect 17596 6776 17606 6862
rect 18032 6776 18042 6862
rect 18110 6776 18120 6862
rect 18550 6776 18560 6862
rect 18628 6776 18638 6862
rect 19066 6776 19076 6862
rect 19144 6776 19154 6862
rect 22378 6402 22578 6602
rect 7900 6270 19098 6320
rect 13376 6212 13592 6270
rect 3708 6146 5226 6204
rect 5588 6146 7106 6204
rect 7900 6162 19098 6212
rect 3708 6104 3766 6146
rect 7045 6104 7103 6146
rect 3708 6046 5226 6104
rect 5594 6046 7112 6104
rect 3708 5788 3766 6046
rect 4018 5954 4028 6014
rect 4092 5954 4102 6014
rect 4254 5954 4264 6014
rect 4328 5954 4338 6014
rect 4490 5954 4500 6014
rect 4564 5954 4574 6014
rect 4726 5954 4736 6014
rect 4800 5954 4810 6014
rect 4962 5954 4972 6014
rect 5036 5954 5046 6014
rect 5198 5954 5208 6014
rect 5272 5954 5282 6014
rect 5526 5956 5536 6014
rect 5600 5956 5610 6014
rect 5762 5956 5772 6014
rect 5836 5956 5846 6014
rect 5998 5956 6008 6014
rect 6072 5956 6082 6014
rect 6234 5956 6244 6014
rect 6308 5956 6318 6014
rect 6468 5956 6478 6014
rect 6542 5956 6552 6014
rect 6706 5956 6716 6014
rect 6780 5956 6790 6014
rect 4134 5824 4144 5884
rect 4214 5824 4224 5884
rect 4370 5824 4380 5884
rect 4450 5824 4460 5884
rect 4606 5824 4616 5884
rect 4686 5824 4696 5884
rect 4842 5824 4852 5884
rect 4922 5824 4932 5884
rect 5078 5824 5088 5884
rect 5158 5824 5168 5884
rect 5646 5826 5656 5886
rect 5716 5826 5726 5886
rect 5882 5826 5892 5886
rect 5952 5826 5962 5886
rect 6118 5826 6128 5886
rect 6188 5826 6198 5886
rect 6356 5826 6366 5886
rect 6426 5826 6436 5886
rect 6590 5826 6600 5886
rect 6660 5826 6670 5886
rect 7045 5788 7103 6046
rect 7834 6026 7844 6112
rect 7912 6026 7922 6112
rect 8350 6026 8360 6112
rect 8428 6026 8438 6112
rect 8866 6026 8876 6112
rect 8944 6026 8954 6112
rect 9382 6026 9392 6112
rect 9460 6026 9470 6112
rect 9898 6026 9908 6112
rect 9976 6026 9986 6112
rect 10414 6026 10424 6112
rect 10492 6026 10502 6112
rect 10928 6026 10938 6112
rect 11006 6026 11016 6112
rect 11446 6026 11456 6112
rect 11524 6026 11534 6112
rect 11962 6026 11972 6112
rect 12040 6026 12050 6112
rect 12478 6026 12488 6112
rect 12556 6026 12566 6112
rect 12996 6026 13006 6112
rect 13074 6026 13084 6112
rect 3708 5730 5226 5788
rect 5588 5730 7106 5788
rect 4537 5684 4807 5693
rect 4537 5626 4556 5684
rect 4794 5626 4807 5684
rect 1110 5338 1218 5538
rect 546 5132 1218 5338
rect 1502 5172 1606 5528
rect 1878 5172 1982 5524
rect 1502 5068 1982 5172
rect 2290 5178 2404 5528
rect 2689 5178 2803 5549
rect 2290 5064 2803 5178
rect 3088 5174 3188 5536
rect 4537 5420 4807 5626
rect 6012 5686 6297 5694
rect 6012 5624 6034 5686
rect 6276 5624 6297 5686
rect 7045 5652 7103 5730
rect 5009 5420 5172 5426
rect 5650 5420 5813 5426
rect 6012 5420 6297 5624
rect 7025 5543 7124 5652
rect 13376 5584 13592 6162
rect 13906 6026 13916 6112
rect 13984 6026 13994 6112
rect 14422 6028 14432 6114
rect 14500 6028 14510 6114
rect 14938 6028 14948 6114
rect 15016 6028 15026 6114
rect 15454 6028 15464 6114
rect 15532 6028 15542 6114
rect 15970 6028 15980 6114
rect 16048 6028 16058 6114
rect 16486 6028 16496 6114
rect 16564 6028 16574 6114
rect 17002 6028 17012 6114
rect 17080 6028 17090 6114
rect 17518 6028 17528 6114
rect 17596 6028 17606 6114
rect 18034 6028 18044 6114
rect 18112 6028 18122 6114
rect 18550 6028 18560 6114
rect 18628 6028 18638 6114
rect 19066 6028 19076 6114
rect 19144 6028 19154 6114
rect 4537 5257 5009 5420
rect 4537 5203 4807 5257
rect 5009 5251 5172 5257
rect 5649 5257 5650 5420
rect 5813 5257 6297 5420
rect 5649 5256 6297 5257
rect 5650 5251 5813 5256
rect 6012 5196 6297 5256
rect 3084 5168 3520 5174
rect 3084 5078 3636 5168
rect 3088 5075 3188 5078
rect 814 5000 3242 5014
rect 814 4998 2258 5000
rect 814 4942 1078 4998
rect 1242 4942 1472 4998
rect 1636 4942 1866 4998
rect 2030 4942 2258 4998
rect 2428 4942 2670 5000
rect 2834 4942 3062 5000
rect 3224 4942 3242 5000
rect 814 4930 3242 4942
rect 98 4358 298 4386
rect 475 4363 645 4369
rect 98 4199 475 4358
rect 98 4186 298 4199
rect 475 4187 645 4193
rect 814 3582 898 4930
rect 3428 4072 3636 5078
rect 3879 4817 4049 4823
rect 6989 4817 7159 5543
rect 7898 5534 19096 5584
rect 13376 5476 13592 5534
rect 7900 5426 19098 5476
rect 7834 5298 7844 5384
rect 7912 5298 7922 5384
rect 8350 5298 8360 5384
rect 8428 5298 8438 5384
rect 8868 5298 8878 5384
rect 8946 5298 8956 5384
rect 9382 5298 9392 5384
rect 9460 5298 9470 5384
rect 9898 5300 9908 5386
rect 9976 5300 9986 5386
rect 10416 5300 10426 5386
rect 10494 5300 10504 5386
rect 10930 5300 10940 5386
rect 11008 5300 11018 5386
rect 11448 5300 11458 5386
rect 11526 5300 11536 5386
rect 11962 5300 11972 5386
rect 12040 5300 12050 5386
rect 12478 5300 12488 5386
rect 12556 5300 12566 5386
rect 12996 5300 13006 5386
rect 13074 5300 13084 5386
rect 13376 4846 13592 5426
rect 13906 5300 13916 5386
rect 13984 5300 13994 5386
rect 14424 5300 14434 5386
rect 14502 5300 14512 5386
rect 14938 5300 14948 5386
rect 15016 5300 15026 5386
rect 15454 5300 15464 5386
rect 15532 5300 15542 5386
rect 15970 5300 15980 5386
rect 16048 5300 16058 5386
rect 16486 5300 16496 5386
rect 16564 5300 16574 5386
rect 17002 5300 17012 5386
rect 17080 5300 17090 5386
rect 17518 5300 17528 5386
rect 17596 5300 17606 5386
rect 18034 5300 18044 5386
rect 18112 5300 18122 5386
rect 18550 5300 18560 5386
rect 18628 5300 18638 5386
rect 19066 5300 19076 5386
rect 19144 5300 19154 5386
rect 4049 4647 7159 4817
rect 7900 4796 19098 4846
rect 3879 4641 4049 4647
rect 1533 4002 1682 4008
rect 3428 4002 6574 4072
rect 1682 3864 6574 4002
rect 1682 3853 3678 3864
rect 1533 3847 1682 3853
rect 1218 3627 6304 3630
rect 6495 3627 6569 3864
rect 49 3556 1148 3582
rect 1218 3556 6569 3627
rect 49 3292 1068 3556
rect 1142 3292 1148 3556
rect 6255 3553 6569 3556
rect 1190 3460 1200 3522
rect 1256 3460 1266 3522
rect 2106 3460 2116 3522
rect 2172 3460 2182 3522
rect 3022 3460 3032 3522
rect 3088 3460 3098 3522
rect 3938 3460 3948 3522
rect 4004 3460 4014 3522
rect 4852 3456 4862 3518
rect 4918 3456 4928 3518
rect 5768 3458 5778 3520
rect 5834 3458 5844 3520
rect 1642 3318 1652 3374
rect 1722 3318 1732 3374
rect 2558 3318 2568 3374
rect 2638 3318 2648 3374
rect 3472 3320 3482 3376
rect 3552 3320 3562 3376
rect 4390 3318 4400 3374
rect 4470 3318 4480 3374
rect 5306 3318 5316 3374
rect 5386 3318 5396 3374
rect 49 3272 1148 3292
rect 6495 3282 6569 3553
rect 6986 3510 7159 4647
rect 7410 4232 7416 4392
rect 7576 4232 7582 4392
rect 7416 3899 7576 4232
rect 13376 4122 13592 4796
rect 22380 4698 22580 4898
rect 7606 3899 10316 3900
rect 7412 3831 10316 3899
rect 6986 3461 7004 3510
rect 49 1528 359 3272
rect 575 3270 768 3272
rect 1222 3208 6569 3282
rect 6983 3374 7004 3461
rect 7140 3374 7159 3510
rect 6983 3356 7159 3374
rect 7606 3830 10316 3831
rect 7606 3370 7676 3830
rect 8036 3706 8046 3790
rect 8106 3706 8116 3790
rect 8272 3706 8282 3790
rect 8342 3706 8352 3790
rect 8506 3706 8516 3790
rect 8576 3706 8586 3790
rect 8742 3706 8752 3790
rect 8812 3706 8822 3790
rect 8978 3706 8988 3790
rect 9048 3706 9058 3790
rect 9214 3706 9224 3790
rect 9284 3706 9294 3790
rect 9450 3706 9460 3790
rect 9520 3706 9530 3790
rect 9686 3706 9696 3790
rect 9756 3706 9766 3790
rect 9922 3706 9932 3790
rect 9992 3706 10002 3790
rect 10158 3706 10168 3790
rect 10228 3706 10238 3790
rect 7912 3402 7922 3486
rect 7990 3402 8000 3486
rect 8148 3402 8158 3486
rect 8226 3402 8236 3486
rect 8386 3402 8396 3486
rect 8464 3402 8474 3486
rect 8622 3402 8632 3486
rect 8700 3402 8710 3486
rect 8858 3402 8868 3486
rect 8936 3402 8946 3486
rect 9094 3402 9104 3486
rect 9172 3402 9182 3486
rect 9330 3402 9340 3486
rect 9408 3402 9418 3486
rect 9566 3404 9576 3488
rect 9644 3404 9654 3488
rect 9802 3404 9812 3488
rect 9880 3404 9890 3488
rect 10038 3404 10048 3488
rect 10116 3404 10126 3488
rect 10274 3404 10284 3488
rect 10352 3404 10362 3488
rect 746 2923 873 2929
rect 746 2664 873 2796
rect 6131 2789 6137 2851
rect 6199 2789 6205 2851
rect 780 2546 838 2664
rect 780 2545 5800 2546
rect 778 2488 5800 2545
rect 778 2230 828 2488
rect 1652 2372 1720 2488
rect 2564 2372 2632 2488
rect 3484 2372 3552 2488
rect 4398 2372 4466 2488
rect 5314 2372 5382 2488
rect 1180 2262 1190 2318
rect 1260 2262 1270 2318
rect 2098 2264 2108 2320
rect 2178 2264 2188 2320
rect 3012 2264 3022 2320
rect 3092 2264 3102 2320
rect 3930 2264 3940 2320
rect 4010 2264 4020 2320
rect 4844 2264 4854 2320
rect 4924 2264 4934 2320
rect 5764 2264 5774 2320
rect 5844 2264 5854 2320
rect 778 2180 5798 2230
rect 1972 2134 2310 2148
rect 1972 2042 2038 2134
rect 2246 2042 2310 2134
rect 575 1528 830 1530
rect 1972 1528 2310 2042
rect 4762 2134 5098 2148
rect 4762 2046 4814 2134
rect 5046 2046 5098 2134
rect 4762 1528 5098 2046
rect 6137 1528 6199 2789
rect 6410 2554 6525 3208
rect 6983 3090 7158 3356
rect 7606 3300 10316 3370
rect 8636 3266 9458 3272
rect 8636 3202 8684 3266
rect 9426 3202 9458 3266
rect 8636 3114 9458 3202
rect 8636 3090 8724 3114
rect 6983 3002 8724 3090
rect 6983 2997 7158 3002
rect 6981 2959 7158 2997
rect 6981 2883 7131 2959
rect 6981 2777 7003 2883
rect 7109 2777 7131 2883
rect 6981 2755 7131 2777
rect 6410 2484 11278 2554
rect 6410 2462 6525 2484
rect 6432 2226 6482 2462
rect 7114 2398 7124 2450
rect 7190 2398 7200 2450
rect 8032 2398 8042 2450
rect 8108 2398 8118 2450
rect 8946 2398 8956 2450
rect 9022 2398 9032 2450
rect 9862 2398 9872 2450
rect 9938 2398 9948 2450
rect 10780 2398 10790 2450
rect 10856 2398 10866 2450
rect 6658 2262 6668 2314
rect 6734 2262 6744 2314
rect 7574 2262 7584 2314
rect 7650 2262 7660 2314
rect 8490 2262 8500 2314
rect 8566 2262 8576 2314
rect 9406 2262 9416 2314
rect 9482 2262 9492 2314
rect 10322 2262 10332 2314
rect 10398 2262 10408 2314
rect 11238 2262 11248 2314
rect 11314 2262 11324 2314
rect 6432 2176 11278 2226
rect 7462 2138 7800 2146
rect 7462 2052 7516 2138
rect 7754 2052 7800 2138
rect 7462 1528 7800 2052
rect 10206 2136 10546 2148
rect 10206 2052 10260 2136
rect 10500 2052 10546 2136
rect 10206 1528 10546 2052
rect 12692 2138 13036 2150
rect 12692 2052 12758 2138
rect 12986 2052 13036 2138
rect 11464 2010 11470 2051
rect 11420 1982 11470 2010
rect 11539 2010 11545 2051
rect 11539 1982 11588 2010
rect 11420 1528 11588 1982
rect 12692 1528 13036 2052
rect 15488 2136 15834 2148
rect 15488 2054 15548 2136
rect 15776 2054 15834 2136
rect 15488 1528 15834 2054
rect 17864 2136 18210 2148
rect 17864 2060 17912 2136
rect 18164 2060 18210 2136
rect 17864 2052 18210 2060
rect 20676 2136 21024 2148
rect 20676 2056 20726 2136
rect 20964 2056 21024 2136
rect 17864 1528 18212 2052
rect 20676 1528 21024 2056
rect 10 1494 22586 1528
rect 10 1404 1000 1494
rect 1240 1404 22586 1494
rect 10 1082 22586 1404
rect 17864 1078 18212 1082
<< via1 >>
rect 546 9930 752 10136
rect 3508 10086 3600 10178
rect 7264 10084 7359 10179
rect 13417 10036 13552 10171
rect 3778 9718 3840 9774
rect 4292 9720 4354 9776
rect 4810 9722 4872 9778
rect 4034 9592 4098 9652
rect 4550 9592 4614 9652
rect 5066 9592 5130 9652
rect 5990 9722 6052 9778
rect 6508 9722 6570 9778
rect 7024 9722 7086 9778
rect 7844 9712 7912 9798
rect 8362 9712 8430 9798
rect 8878 9712 8946 9798
rect 9394 9712 9462 9798
rect 9910 9712 9978 9798
rect 10426 9712 10494 9798
rect 10942 9712 11010 9798
rect 11458 9712 11526 9798
rect 11972 9712 12040 9798
rect 12490 9712 12558 9798
rect 13006 9712 13074 9798
rect 5275 9586 5329 9640
rect 5734 9584 5798 9644
rect 6248 9584 6312 9644
rect 6766 9584 6830 9644
rect 13918 9712 13986 9798
rect 14432 9712 14500 9798
rect 14948 9712 15016 9798
rect 15464 9712 15532 9798
rect 15982 9712 16050 9798
rect 16496 9712 16564 9798
rect 17014 9712 17082 9798
rect 17528 9712 17596 9798
rect 18046 9712 18114 9798
rect 18560 9712 18628 9798
rect 19078 9712 19146 9798
rect 7844 8974 7912 9060
rect 8360 8974 8428 9060
rect 8878 8974 8946 9060
rect 9392 8974 9460 9060
rect 9908 8974 9976 9060
rect 10424 8974 10492 9060
rect 10940 8974 11008 9060
rect 11456 8976 11524 9062
rect 11972 8976 12040 9062
rect 12488 8976 12556 9062
rect 13006 8976 13074 9062
rect 13918 8976 13986 9062
rect 14432 8976 14500 9062
rect 14948 8976 15016 9062
rect 15466 8976 15534 9062
rect 15978 8976 16046 9062
rect 16496 8972 16564 9058
rect 17012 8972 17080 9058
rect 17526 8972 17594 9058
rect 18044 8972 18112 9058
rect 18562 8972 18630 9058
rect 19078 8972 19146 9058
rect 7844 8246 7912 8332
rect 8360 8246 8428 8332
rect 8876 8246 8944 8332
rect 9392 8246 9460 8332
rect 9908 8246 9976 8332
rect 10424 8246 10492 8332
rect 10940 8246 11008 8332
rect 11456 8246 11524 8332
rect 11972 8246 12040 8332
rect 12488 8246 12556 8332
rect 13004 8246 13072 8332
rect 546 6937 752 7143
rect 13918 8244 13986 8330
rect 14430 8244 14498 8330
rect 14948 8244 15016 8330
rect 15464 8244 15532 8330
rect 15980 8244 16048 8330
rect 16496 8244 16564 8330
rect 17012 8244 17080 8330
rect 17528 8244 17596 8330
rect 18044 8244 18112 8330
rect 18560 8244 18628 8330
rect 19076 8244 19144 8330
rect 4030 7626 4094 7686
rect 4264 7626 4328 7686
rect 4500 7626 4564 7686
rect 4736 7626 4800 7686
rect 4972 7626 5036 7686
rect 5208 7626 5272 7686
rect 5536 7626 5600 7684
rect 5772 7626 5836 7684
rect 6008 7626 6072 7684
rect 6244 7626 6308 7684
rect 6480 7626 6544 7684
rect 6716 7626 6780 7684
rect 4144 7490 4214 7550
rect 4380 7492 4450 7552
rect 4616 7492 4686 7552
rect 4850 7492 4920 7552
rect 5088 7492 5158 7552
rect 5656 7492 5716 7552
rect 5892 7492 5952 7552
rect 6128 7492 6188 7552
rect 6364 7492 6424 7552
rect 6600 7492 6660 7552
rect 7844 7504 7912 7590
rect 8360 7504 8428 7590
rect 8876 7504 8944 7590
rect 9392 7504 9460 7590
rect 9908 7504 9976 7590
rect 10424 7504 10492 7590
rect 10940 7504 11008 7590
rect 11456 7504 11524 7590
rect 11974 7504 12042 7590
rect 12490 7504 12558 7590
rect 13006 7504 13074 7590
rect 4028 7208 4092 7268
rect 4264 7208 4328 7268
rect 4500 7208 4564 7268
rect 4736 7208 4800 7268
rect 4972 7208 5036 7268
rect 5210 7208 5274 7268
rect 5536 7208 5600 7266
rect 5772 7208 5836 7266
rect 6008 7208 6072 7266
rect 6244 7208 6308 7266
rect 6480 7208 6544 7266
rect 6716 7208 6780 7266
rect 4142 7076 4212 7136
rect 4380 7076 4450 7136
rect 4616 7076 4686 7136
rect 4852 7076 4922 7136
rect 5088 7076 5158 7136
rect 5656 7072 5716 7132
rect 5892 7072 5952 7132
rect 6128 7072 6188 7132
rect 6364 7072 6424 7132
rect 6600 7072 6660 7132
rect 13916 7504 13984 7590
rect 14432 7504 14500 7590
rect 14948 7504 15016 7590
rect 15464 7504 15532 7590
rect 15980 7504 16048 7590
rect 16496 7504 16564 7590
rect 17012 7504 17080 7590
rect 17528 7504 17596 7590
rect 18044 7504 18112 7590
rect 18560 7504 18628 7590
rect 19078 7504 19146 7590
rect 4028 6788 4092 6848
rect 4264 6790 4328 6850
rect 4502 6790 4566 6850
rect 4736 6790 4800 6850
rect 4972 6790 5036 6850
rect 5208 6790 5272 6850
rect 5536 6792 5600 6850
rect 5772 6792 5836 6850
rect 6010 6792 6074 6850
rect 6244 6792 6308 6850
rect 6480 6792 6544 6850
rect 6716 6794 6780 6852
rect 4142 6656 4212 6716
rect 4380 6656 4450 6716
rect 4616 6656 4686 6716
rect 4852 6656 4922 6716
rect 5090 6656 5160 6716
rect 5656 6660 5716 6720
rect 5892 6660 5952 6720
rect 6128 6660 6188 6720
rect 6364 6660 6424 6720
rect 6600 6660 6660 6720
rect 7844 6776 7912 6862
rect 8360 6776 8428 6862
rect 8874 6776 8942 6862
rect 9392 6776 9460 6862
rect 9908 6776 9976 6862
rect 10424 6776 10492 6862
rect 10940 6776 11008 6862
rect 11456 6776 11524 6862
rect 11972 6776 12040 6862
rect 12488 6776 12556 6862
rect 13006 6776 13074 6862
rect 4028 6374 4092 6434
rect 4264 6374 4328 6434
rect 4500 6374 4564 6434
rect 4736 6374 4800 6434
rect 4972 6374 5036 6434
rect 5208 6374 5272 6434
rect 5536 6376 5600 6434
rect 5772 6376 5836 6434
rect 6008 6376 6072 6434
rect 6244 6376 6308 6434
rect 6480 6376 6544 6434
rect 6716 6376 6780 6434
rect 4144 6240 4214 6300
rect 4380 6240 4450 6300
rect 4616 6240 4686 6300
rect 4852 6240 4922 6300
rect 5088 6240 5158 6300
rect 5656 6244 5716 6304
rect 5892 6244 5952 6304
rect 6128 6244 6188 6304
rect 6364 6244 6424 6304
rect 6600 6244 6660 6304
rect 13916 6776 13984 6862
rect 14430 6776 14498 6862
rect 14948 6776 15016 6862
rect 15464 6776 15532 6862
rect 15980 6776 16048 6862
rect 16498 6776 16566 6862
rect 17010 6776 17078 6862
rect 17528 6776 17596 6862
rect 18042 6776 18110 6862
rect 18560 6776 18628 6862
rect 19076 6776 19144 6862
rect 4028 5954 4092 6014
rect 4264 5954 4328 6014
rect 4500 5954 4564 6014
rect 4736 5954 4800 6014
rect 4972 5954 5036 6014
rect 5208 5954 5272 6014
rect 5536 5956 5600 6014
rect 5772 5956 5836 6014
rect 6008 5956 6072 6014
rect 6244 5956 6308 6014
rect 6478 5956 6542 6014
rect 6716 5956 6780 6014
rect 4144 5824 4214 5884
rect 4380 5824 4450 5884
rect 4616 5824 4686 5884
rect 4852 5824 4922 5884
rect 5088 5824 5158 5884
rect 5656 5826 5716 5886
rect 5892 5826 5952 5886
rect 6128 5826 6188 5886
rect 6366 5826 6426 5886
rect 6600 5826 6660 5886
rect 7844 6026 7912 6112
rect 8360 6026 8428 6112
rect 8876 6026 8944 6112
rect 9392 6026 9460 6112
rect 9908 6026 9976 6112
rect 10424 6026 10492 6112
rect 10938 6026 11006 6112
rect 11456 6026 11524 6112
rect 11972 6026 12040 6112
rect 12488 6026 12556 6112
rect 13006 6026 13074 6112
rect 13916 6026 13984 6112
rect 14432 6028 14500 6114
rect 14948 6028 15016 6114
rect 15464 6028 15532 6114
rect 15980 6028 16048 6114
rect 16496 6028 16564 6114
rect 17012 6028 17080 6114
rect 17528 6028 17596 6114
rect 18044 6028 18112 6114
rect 18560 6028 18628 6114
rect 19076 6028 19144 6114
rect 5009 5257 5172 5420
rect 5650 5257 5813 5420
rect 475 4193 645 4363
rect 7844 5298 7912 5384
rect 8360 5298 8428 5384
rect 8878 5298 8946 5384
rect 9392 5298 9460 5384
rect 9908 5300 9976 5386
rect 10426 5300 10494 5386
rect 10940 5300 11008 5386
rect 11458 5300 11526 5386
rect 11972 5300 12040 5386
rect 12488 5300 12556 5386
rect 13006 5300 13074 5386
rect 13916 5300 13984 5386
rect 14434 5300 14502 5386
rect 14948 5300 15016 5386
rect 15464 5300 15532 5386
rect 15980 5300 16048 5386
rect 16496 5300 16564 5386
rect 17012 5300 17080 5386
rect 17528 5300 17596 5386
rect 18044 5300 18112 5386
rect 18560 5300 18628 5386
rect 19076 5300 19144 5386
rect 3879 4647 4049 4817
rect 1533 3853 1682 4002
rect 1200 3460 1256 3522
rect 2116 3460 2172 3522
rect 3032 3460 3088 3522
rect 3948 3460 4004 3522
rect 4862 3456 4918 3518
rect 5778 3458 5834 3520
rect 1652 3318 1722 3374
rect 2568 3318 2638 3374
rect 3482 3320 3552 3376
rect 4400 3318 4470 3374
rect 5316 3318 5386 3374
rect 7416 4232 7576 4392
rect 7004 3374 7140 3510
rect 8046 3706 8106 3790
rect 8282 3706 8342 3790
rect 8516 3706 8576 3790
rect 8752 3706 8812 3790
rect 8988 3706 9048 3790
rect 9224 3706 9284 3790
rect 9460 3706 9520 3790
rect 9696 3706 9756 3790
rect 9932 3706 9992 3790
rect 10168 3706 10228 3790
rect 7922 3402 7990 3486
rect 8158 3402 8226 3486
rect 8396 3402 8464 3486
rect 8632 3402 8700 3486
rect 8868 3402 8936 3486
rect 9104 3402 9172 3486
rect 9340 3402 9408 3486
rect 9576 3404 9644 3488
rect 9812 3404 9880 3488
rect 10048 3404 10116 3488
rect 10284 3404 10352 3488
rect 746 2796 873 2923
rect 6137 2789 6199 2851
rect 1190 2262 1260 2318
rect 2108 2264 2178 2320
rect 3022 2264 3092 2320
rect 3940 2264 4010 2320
rect 4854 2264 4924 2320
rect 5774 2264 5844 2320
rect 7003 2777 7109 2883
rect 7124 2398 7190 2450
rect 8042 2398 8108 2450
rect 8956 2398 9022 2450
rect 9872 2398 9938 2450
rect 10790 2398 10856 2450
rect 6668 2262 6734 2314
rect 7584 2262 7650 2314
rect 8500 2262 8566 2314
rect 9416 2262 9482 2314
rect 10332 2262 10398 2314
rect 11248 2262 11314 2314
rect 11470 1982 11539 2051
rect 1000 1404 1240 1494
<< metal2 >>
rect 3508 10178 3600 10184
rect 540 9930 546 10136
rect 752 9930 758 10136
rect 546 7143 752 9930
rect 3508 9800 3600 10086
rect 7264 10179 7359 10185
rect 7264 9802 7359 10084
rect 13417 10171 13552 10177
rect 3508 9782 3662 9800
rect 3778 9782 3840 9784
rect 4292 9782 4354 9786
rect 4810 9782 4872 9788
rect 5990 9782 6052 9788
rect 6508 9782 6570 9788
rect 7024 9782 7086 9788
rect 7197 9782 7359 9802
rect 3508 9778 5136 9782
rect 3508 9776 4810 9778
rect 3508 9774 4292 9776
rect 3508 9726 3778 9774
rect 3508 9708 3662 9726
rect 3840 9726 4292 9774
rect 3778 9708 3840 9718
rect 4354 9726 4810 9776
rect 4292 9710 4354 9720
rect 4872 9726 5136 9778
rect 5724 9778 7359 9782
rect 5724 9726 5990 9778
rect 4810 9712 4872 9722
rect 6052 9726 6508 9778
rect 5990 9712 6052 9722
rect 6570 9726 7024 9778
rect 6508 9712 6570 9722
rect 7086 9726 7359 9778
rect 7024 9712 7086 9722
rect 7197 9707 7359 9726
rect 7844 9798 7912 9808
rect 8362 9798 8430 9808
rect 8878 9798 8946 9808
rect 9394 9798 9462 9808
rect 9910 9798 9978 9808
rect 10426 9798 10494 9808
rect 10942 9798 11010 9808
rect 11458 9798 11526 9808
rect 11972 9798 12040 9808
rect 12490 9798 12558 9808
rect 13006 9798 13074 9808
rect 13417 9798 13552 10036
rect 13918 9798 13986 9808
rect 14432 9798 14500 9808
rect 14948 9798 15016 9808
rect 15464 9798 15532 9808
rect 15982 9798 16050 9808
rect 16496 9798 16564 9808
rect 17014 9798 17082 9808
rect 17528 9798 17596 9808
rect 18046 9798 18114 9808
rect 18560 9798 18628 9808
rect 19078 9798 19146 9808
rect 7912 9722 8362 9798
rect 7844 9702 7912 9712
rect 8430 9722 8878 9798
rect 8362 9702 8430 9712
rect 8946 9722 9394 9798
rect 8878 9702 8946 9712
rect 9462 9722 9910 9798
rect 9394 9702 9462 9712
rect 9978 9722 10426 9798
rect 9910 9702 9978 9712
rect 10494 9722 10942 9798
rect 10426 9702 10494 9712
rect 11010 9722 11458 9798
rect 10942 9702 11010 9712
rect 11526 9722 11972 9798
rect 11458 9702 11526 9712
rect 12040 9722 12490 9798
rect 11972 9702 12040 9712
rect 12558 9722 13006 9798
rect 12490 9702 12558 9712
rect 13074 9722 13918 9798
rect 13006 9702 13074 9712
rect 4034 9652 4098 9662
rect 3505 9640 3567 9644
rect 3505 9592 4034 9640
rect 4550 9652 4614 9662
rect 4098 9592 4550 9640
rect 5066 9652 5130 9662
rect 4614 9592 5066 9640
rect 5734 9644 5798 9654
rect 5130 9592 5275 9640
rect 3505 9586 5275 9592
rect 5329 9586 5335 9640
rect 3505 9375 3567 9586
rect 4034 9582 4098 9586
rect 4550 9582 4614 9586
rect 5066 9582 5130 9586
rect 5722 9584 5734 9632
rect 6248 9644 6312 9654
rect 5798 9584 6248 9632
rect 6766 9644 6830 9654
rect 6312 9584 6766 9632
rect 6830 9584 7349 9632
rect 5722 9578 7349 9584
rect 5734 9574 5798 9578
rect 6248 9574 6312 9578
rect 6766 9574 6830 9578
rect 7295 9421 7349 9578
rect 3465 8905 3607 9375
rect 7249 8921 7395 9421
rect 7844 9060 7912 9070
rect 8360 9060 8428 9070
rect 8878 9060 8946 9070
rect 9392 9060 9460 9070
rect 9908 9060 9976 9070
rect 10424 9060 10492 9070
rect 10940 9060 11008 9070
rect 11456 9062 11524 9072
rect 7912 8984 8360 9060
rect 7844 8964 7912 8974
rect 8428 8984 8878 9060
rect 8360 8964 8428 8974
rect 8946 8984 9392 9060
rect 8878 8964 8946 8974
rect 9460 8984 9908 9060
rect 9392 8964 9460 8974
rect 9976 8984 10424 9060
rect 9908 8964 9976 8974
rect 10492 8984 10940 9060
rect 10424 8964 10492 8974
rect 11008 8984 11456 9060
rect 10940 8964 11008 8974
rect 11972 9062 12040 9072
rect 11524 8984 11972 9060
rect 11456 8966 11524 8976
rect 12488 9062 12556 9072
rect 12040 8984 12488 9060
rect 11972 8966 12040 8976
rect 13006 9062 13074 9072
rect 12556 8984 13006 9060
rect 12488 8966 12556 8976
rect 13242 9060 13318 9722
rect 13417 9693 13552 9722
rect 13657 9060 13731 9722
rect 13986 9722 14432 9798
rect 13918 9702 13986 9712
rect 14500 9722 14948 9798
rect 14432 9702 14500 9712
rect 15016 9722 15464 9798
rect 14948 9702 15016 9712
rect 15532 9722 15982 9798
rect 15464 9702 15532 9712
rect 16050 9722 16496 9798
rect 15982 9702 16050 9712
rect 16564 9722 17014 9798
rect 16496 9702 16564 9712
rect 17082 9722 17528 9798
rect 17014 9702 17082 9712
rect 17596 9722 18046 9798
rect 17528 9702 17596 9712
rect 18114 9722 18560 9798
rect 18046 9702 18114 9712
rect 18628 9722 19078 9798
rect 18560 9702 18628 9712
rect 19146 9722 19158 9798
rect 19078 9702 19146 9712
rect 13918 9062 13986 9072
rect 13074 8984 13918 9060
rect 13006 8966 13074 8976
rect 3465 8763 3771 8905
rect 3629 7694 3771 8763
rect 7057 8775 7395 8921
rect 4030 7694 4094 7696
rect 4264 7694 4328 7696
rect 4500 7694 4564 7696
rect 4736 7694 4800 7696
rect 4972 7694 5036 7696
rect 5208 7694 5272 7696
rect 7057 7694 7203 8775
rect 7844 8332 7912 8342
rect 8360 8332 8428 8342
rect 8876 8332 8944 8342
rect 9392 8332 9460 8342
rect 9908 8332 9976 8342
rect 10424 8332 10492 8342
rect 10940 8332 11008 8342
rect 11456 8332 11524 8342
rect 11972 8332 12040 8342
rect 12488 8332 12556 8342
rect 13004 8332 13072 8342
rect 13242 8332 13318 8984
rect 13657 8332 13731 8984
rect 14432 9062 14500 9072
rect 13986 8984 14432 9060
rect 13918 8966 13986 8976
rect 14948 9062 15016 9072
rect 14500 8984 14948 9060
rect 14432 8966 14500 8976
rect 15466 9062 15534 9072
rect 15016 8984 15466 9060
rect 14948 8966 15016 8976
rect 15978 9062 16046 9072
rect 15534 8984 15978 9060
rect 15466 8966 15534 8976
rect 16496 9060 16564 9068
rect 17012 9060 17080 9068
rect 17526 9060 17594 9068
rect 18044 9060 18112 9068
rect 18562 9060 18630 9068
rect 19078 9060 19146 9068
rect 16046 9058 19160 9060
rect 16046 8984 16496 9058
rect 15978 8966 16046 8976
rect 16564 8984 17012 9058
rect 16496 8962 16564 8972
rect 17080 8984 17526 9058
rect 17012 8962 17080 8972
rect 17594 8984 18044 9058
rect 17526 8962 17594 8972
rect 18112 8984 18562 9058
rect 18044 8962 18112 8972
rect 18630 8984 19078 9058
rect 18562 8962 18630 8972
rect 19146 8984 19160 9058
rect 19078 8962 19146 8972
rect 13918 8332 13986 8340
rect 14430 8332 14498 8340
rect 14948 8332 15016 8340
rect 15464 8332 15532 8340
rect 15980 8332 16048 8340
rect 16496 8332 16564 8340
rect 17012 8332 17080 8340
rect 17528 8332 17596 8340
rect 18044 8332 18112 8340
rect 18560 8332 18628 8340
rect 19076 8332 19144 8340
rect 7912 8256 8360 8332
rect 7844 8236 7912 8246
rect 8428 8256 8876 8332
rect 8360 8236 8428 8246
rect 8944 8256 9392 8332
rect 8876 8236 8944 8246
rect 9460 8256 9908 8332
rect 9392 8236 9460 8246
rect 9976 8256 10424 8332
rect 9908 8236 9976 8246
rect 10492 8256 10940 8332
rect 10424 8236 10492 8246
rect 11008 8256 11456 8332
rect 10940 8236 11008 8246
rect 11524 8256 11972 8332
rect 11456 8236 11524 8246
rect 12040 8256 12488 8332
rect 11972 8236 12040 8246
rect 12556 8256 13004 8332
rect 12488 8236 12556 8246
rect 13072 8330 19160 8332
rect 13072 8256 13918 8330
rect 13004 8236 13072 8246
rect 546 6931 752 6937
rect 3615 7686 5278 7694
rect 3615 7636 4030 7686
rect 3615 7274 3673 7636
rect 4094 7636 4264 7686
rect 4030 7616 4094 7626
rect 4328 7636 4500 7686
rect 4264 7616 4328 7626
rect 4564 7636 4736 7686
rect 4500 7616 4564 7626
rect 4800 7636 4972 7686
rect 4736 7616 4800 7626
rect 5036 7636 5208 7686
rect 4972 7616 5036 7626
rect 5272 7636 5278 7686
rect 5524 7684 7216 7694
rect 5524 7638 5536 7684
rect 5208 7616 5272 7626
rect 5600 7638 5772 7684
rect 5536 7616 5600 7626
rect 5836 7638 6008 7684
rect 5772 7616 5836 7626
rect 6072 7638 6244 7684
rect 6008 7616 6072 7626
rect 6308 7638 6480 7684
rect 6244 7616 6308 7626
rect 6544 7638 6716 7684
rect 6480 7616 6544 7626
rect 6780 7638 7216 7684
rect 6716 7616 6780 7626
rect 3836 7547 3918 7560
rect 3836 7487 3847 7547
rect 3907 7546 3918 7547
rect 4144 7550 4214 7560
rect 3907 7490 4144 7546
rect 4380 7552 4450 7562
rect 4214 7492 4380 7546
rect 4616 7552 4686 7562
rect 4450 7492 4616 7546
rect 4850 7552 4920 7562
rect 4686 7492 4850 7546
rect 5088 7552 5158 7562
rect 4920 7492 5088 7546
rect 5656 7552 5716 7562
rect 5158 7544 5278 7546
rect 5375 7544 5446 7550
rect 5158 7540 5532 7544
rect 5158 7492 5656 7540
rect 5892 7552 5952 7562
rect 5716 7492 5892 7540
rect 6128 7552 6188 7562
rect 5952 7492 6128 7540
rect 6364 7552 6424 7562
rect 6188 7492 6364 7540
rect 6600 7552 6660 7562
rect 6424 7492 6600 7540
rect 6901 7540 6910 7542
rect 6660 7492 6910 7540
rect 4214 7490 6910 7492
rect 3907 7488 6910 7490
rect 3907 7487 3918 7488
rect 3836 7476 3918 7487
rect 4144 7480 4214 7488
rect 4380 7482 4450 7488
rect 4616 7482 4686 7488
rect 4850 7482 4920 7488
rect 5088 7482 5158 7488
rect 5272 7484 6910 7488
rect 4028 7274 4092 7278
rect 4264 7274 4328 7278
rect 4500 7274 4564 7278
rect 4736 7274 4800 7278
rect 4972 7274 5036 7278
rect 5210 7274 5274 7278
rect 3615 7268 5278 7274
rect 3615 7216 4028 7268
rect 3615 6854 3673 7216
rect 4092 7216 4264 7268
rect 4028 7198 4092 7208
rect 4328 7216 4500 7268
rect 4264 7198 4328 7208
rect 4564 7216 4736 7268
rect 4500 7198 4564 7208
rect 4800 7216 4972 7268
rect 4736 7198 4800 7208
rect 5036 7216 5210 7268
rect 4972 7198 5036 7208
rect 5274 7216 5278 7268
rect 5210 7198 5274 7208
rect 3836 7129 3918 7144
rect 3836 7069 3847 7129
rect 3907 7128 3918 7129
rect 4142 7136 4212 7146
rect 3907 7076 4142 7128
rect 4380 7136 4450 7146
rect 4212 7076 4380 7128
rect 4616 7136 4686 7146
rect 4450 7076 4616 7128
rect 4852 7136 4922 7146
rect 4686 7076 4852 7128
rect 5088 7136 5158 7146
rect 4922 7076 5088 7128
rect 5375 7128 5446 7484
rect 5656 7482 5716 7484
rect 5892 7482 5952 7484
rect 6128 7482 6188 7484
rect 6364 7482 6424 7484
rect 6600 7482 6660 7484
rect 6901 7482 6910 7484
rect 6970 7482 6979 7542
rect 7155 7276 7210 7638
rect 7844 7590 7912 7600
rect 8360 7590 8428 7600
rect 8876 7590 8944 7600
rect 9392 7590 9460 7600
rect 9908 7590 9976 7600
rect 10424 7590 10492 7600
rect 10940 7590 11008 7600
rect 11456 7590 11524 7600
rect 11974 7590 12042 7600
rect 12490 7590 12558 7600
rect 13006 7590 13074 7600
rect 13242 7590 13318 8256
rect 13657 7590 13731 8256
rect 13986 8256 14430 8330
rect 13918 8234 13986 8244
rect 14498 8256 14948 8330
rect 14430 8234 14498 8244
rect 15016 8256 15464 8330
rect 14948 8234 15016 8244
rect 15532 8256 15980 8330
rect 15464 8234 15532 8244
rect 16048 8256 16496 8330
rect 15980 8234 16048 8244
rect 16564 8256 17012 8330
rect 16496 8234 16564 8244
rect 17080 8256 17528 8330
rect 17012 8234 17080 8244
rect 17596 8256 18044 8330
rect 17528 8234 17596 8244
rect 18112 8256 18560 8330
rect 18044 8234 18112 8244
rect 18628 8256 19076 8330
rect 18560 8234 18628 8244
rect 19144 8256 19160 8330
rect 19076 8234 19144 8244
rect 13916 7590 13984 7600
rect 14432 7590 14500 7600
rect 14948 7590 15016 7600
rect 15464 7590 15532 7600
rect 15980 7590 16048 7600
rect 16496 7590 16564 7600
rect 17012 7590 17080 7600
rect 17528 7590 17596 7600
rect 18044 7590 18112 7600
rect 18560 7590 18628 7600
rect 19078 7590 19146 7600
rect 7912 7514 8360 7590
rect 7844 7494 7912 7504
rect 8428 7514 8876 7590
rect 8360 7494 8428 7504
rect 8944 7514 9392 7590
rect 8876 7494 8944 7504
rect 9460 7514 9908 7590
rect 9392 7494 9460 7504
rect 9976 7514 10424 7590
rect 9908 7494 9976 7504
rect 10492 7514 10940 7590
rect 10424 7494 10492 7504
rect 11008 7514 11456 7590
rect 10940 7494 11008 7504
rect 11524 7514 11974 7590
rect 11456 7494 11524 7504
rect 12042 7514 12490 7590
rect 11974 7494 12042 7504
rect 12558 7514 13006 7590
rect 12490 7494 12558 7504
rect 13074 7514 13916 7590
rect 13006 7494 13074 7504
rect 5524 7266 7210 7276
rect 5524 7220 5536 7266
rect 5600 7220 5772 7266
rect 5536 7198 5600 7208
rect 5836 7220 6008 7266
rect 5772 7198 5836 7208
rect 6072 7220 6244 7266
rect 6008 7198 6072 7208
rect 6308 7220 6480 7266
rect 6244 7198 6308 7208
rect 6544 7220 6716 7266
rect 6480 7198 6544 7208
rect 6780 7220 7210 7266
rect 6716 7198 6780 7208
rect 5656 7132 5716 7142
rect 5158 7122 5532 7128
rect 5158 7076 5656 7122
rect 3907 7072 5656 7076
rect 5892 7132 5952 7142
rect 5716 7072 5892 7122
rect 6128 7132 6188 7142
rect 5952 7072 6128 7122
rect 6364 7132 6424 7142
rect 6188 7072 6364 7122
rect 6600 7132 6660 7142
rect 6424 7072 6600 7122
rect 6898 7124 6980 7136
rect 6898 7122 6910 7124
rect 6660 7072 6910 7122
rect 3907 7070 6910 7072
rect 3907 7069 3918 7070
rect 3836 7060 3918 7069
rect 4142 7066 4212 7070
rect 4380 7066 4450 7070
rect 4616 7066 4686 7070
rect 4852 7066 4922 7070
rect 5088 7066 5158 7070
rect 5274 7066 6910 7070
rect 4028 6854 4092 6858
rect 4264 6854 4328 6860
rect 4502 6854 4566 6860
rect 4736 6854 4800 6860
rect 4972 6854 5036 6860
rect 5208 6854 5272 6860
rect 3615 6850 5278 6854
rect 3615 6848 4264 6850
rect 3615 6796 4028 6848
rect 3615 6440 3673 6796
rect 4092 6796 4264 6848
rect 4028 6778 4092 6788
rect 4328 6796 4502 6850
rect 4264 6780 4328 6790
rect 4566 6796 4736 6850
rect 4502 6780 4566 6790
rect 4800 6796 4972 6850
rect 4736 6780 4800 6790
rect 5036 6796 5208 6850
rect 4972 6780 5036 6790
rect 5272 6796 5278 6850
rect 5208 6780 5272 6790
rect 3836 6709 3918 6720
rect 3836 6649 3847 6709
rect 3907 6708 3918 6709
rect 4142 6716 4212 6726
rect 3907 6656 4142 6708
rect 4380 6716 4450 6726
rect 4212 6656 4380 6708
rect 4616 6716 4686 6726
rect 4450 6656 4616 6708
rect 4852 6716 4922 6726
rect 4686 6656 4852 6708
rect 5090 6716 5160 6726
rect 4922 6656 5090 6708
rect 5375 6708 5446 7066
rect 5656 7062 5716 7066
rect 5892 7062 5952 7066
rect 6128 7062 6188 7066
rect 6364 7062 6424 7066
rect 6600 7062 6660 7066
rect 6898 7064 6910 7066
rect 6970 7064 6980 7124
rect 6898 7054 6980 7064
rect 5536 6858 5600 6860
rect 5772 6858 5836 6860
rect 6010 6858 6074 6860
rect 6244 6858 6308 6860
rect 6480 6858 6544 6860
rect 6716 6858 6780 6862
rect 7155 6858 7210 7220
rect 5524 6852 7210 6858
rect 5524 6850 6716 6852
rect 5524 6802 5536 6850
rect 5600 6802 5772 6850
rect 5536 6782 5600 6792
rect 5836 6802 6010 6850
rect 5772 6782 5836 6792
rect 6074 6802 6244 6850
rect 6010 6782 6074 6792
rect 6308 6802 6480 6850
rect 6244 6782 6308 6792
rect 6544 6802 6716 6850
rect 6480 6782 6544 6792
rect 6780 6802 7210 6852
rect 6716 6784 6780 6794
rect 5656 6720 5716 6730
rect 5524 6708 5656 6710
rect 5160 6660 5656 6708
rect 5892 6720 5952 6730
rect 5716 6660 5892 6710
rect 6128 6720 6188 6730
rect 5952 6660 6128 6710
rect 6364 6720 6424 6730
rect 6188 6660 6364 6710
rect 6600 6720 6660 6730
rect 6424 6660 6600 6710
rect 6898 6712 6980 6722
rect 6898 6710 6910 6712
rect 6660 6660 6910 6710
rect 5160 6656 6910 6660
rect 3907 6654 6910 6656
rect 3907 6650 5278 6654
rect 3907 6649 3918 6650
rect 3836 6636 3918 6649
rect 4142 6646 4212 6650
rect 4380 6646 4450 6650
rect 4616 6646 4686 6650
rect 4852 6646 4922 6650
rect 5090 6646 5160 6650
rect 4028 6440 4092 6444
rect 4264 6440 4328 6444
rect 4500 6440 4564 6444
rect 4736 6440 4800 6444
rect 4972 6440 5036 6444
rect 5208 6440 5272 6444
rect 3615 6434 5278 6440
rect 3615 6382 4028 6434
rect 3615 6023 3673 6382
rect 4092 6382 4264 6434
rect 4028 6364 4092 6374
rect 4328 6382 4500 6434
rect 4264 6364 4328 6374
rect 4564 6382 4736 6434
rect 4500 6364 4564 6374
rect 4800 6382 4972 6434
rect 4736 6364 4800 6374
rect 5036 6382 5208 6434
rect 4972 6364 5036 6374
rect 5272 6382 5278 6434
rect 5208 6364 5272 6374
rect 3836 6291 3918 6304
rect 3836 6231 3847 6291
rect 3907 6290 3918 6291
rect 4144 6300 4214 6310
rect 3907 6240 4144 6290
rect 4380 6300 4450 6310
rect 4214 6240 4380 6290
rect 4616 6300 4686 6310
rect 4450 6240 4616 6290
rect 4852 6300 4922 6310
rect 4686 6240 4852 6290
rect 5088 6300 5158 6310
rect 4922 6240 5088 6290
rect 5375 6290 5446 6654
rect 5656 6650 5716 6654
rect 5892 6650 5952 6654
rect 6128 6650 6188 6654
rect 6364 6650 6424 6654
rect 6600 6650 6660 6654
rect 6898 6652 6910 6654
rect 6970 6652 6980 6712
rect 6898 6640 6980 6652
rect 5536 6440 5600 6444
rect 5772 6440 5836 6444
rect 6008 6440 6072 6444
rect 6244 6440 6308 6444
rect 6480 6440 6544 6444
rect 6716 6440 6780 6444
rect 7155 6440 7210 6802
rect 7844 6862 7912 6872
rect 8360 6862 8428 6872
rect 8874 6862 8942 6872
rect 9392 6862 9460 6872
rect 9908 6862 9976 6872
rect 10424 6862 10492 6872
rect 10940 6862 11008 6872
rect 11456 6862 11524 6872
rect 11972 6862 12040 6872
rect 12488 6862 12556 6872
rect 13006 6862 13074 6872
rect 13242 6862 13318 7514
rect 13657 6862 13731 7514
rect 13984 7514 14432 7590
rect 13916 7494 13984 7504
rect 14500 7514 14948 7590
rect 14432 7494 14500 7504
rect 15016 7514 15464 7590
rect 14948 7494 15016 7504
rect 15532 7514 15980 7590
rect 15464 7494 15532 7504
rect 16048 7514 16496 7590
rect 15980 7494 16048 7504
rect 16564 7514 17012 7590
rect 16496 7494 16564 7504
rect 17080 7514 17528 7590
rect 17012 7494 17080 7504
rect 17596 7514 18044 7590
rect 17528 7494 17596 7504
rect 18112 7514 18560 7590
rect 18044 7494 18112 7504
rect 18628 7514 19078 7590
rect 18560 7494 18628 7504
rect 19146 7514 19160 7590
rect 19078 7494 19146 7504
rect 13916 6862 13984 6872
rect 14430 6862 14498 6872
rect 14948 6862 15016 6872
rect 15464 6862 15532 6872
rect 15980 6862 16048 6872
rect 16498 6862 16566 6872
rect 17010 6862 17078 6872
rect 17528 6862 17596 6872
rect 18042 6862 18110 6872
rect 18560 6862 18628 6872
rect 19076 6862 19144 6872
rect 7912 6786 8360 6862
rect 7844 6766 7912 6776
rect 8428 6786 8874 6862
rect 8360 6766 8428 6776
rect 8942 6786 9392 6862
rect 8874 6766 8942 6776
rect 9460 6786 9908 6862
rect 9392 6766 9460 6776
rect 9976 6786 10424 6862
rect 9908 6766 9976 6776
rect 10492 6786 10940 6862
rect 10424 6766 10492 6776
rect 11008 6786 11456 6862
rect 10940 6766 11008 6776
rect 11524 6786 11972 6862
rect 11456 6766 11524 6776
rect 12040 6786 12488 6862
rect 11972 6766 12040 6776
rect 12556 6786 13006 6862
rect 12488 6766 12556 6776
rect 13074 6786 13916 6862
rect 13006 6766 13074 6776
rect 5524 6434 7210 6440
rect 5524 6384 5536 6434
rect 5600 6384 5772 6434
rect 5536 6366 5600 6376
rect 5836 6384 6008 6434
rect 5772 6366 5836 6376
rect 6072 6384 6244 6434
rect 6008 6366 6072 6376
rect 6308 6384 6480 6434
rect 6244 6366 6308 6376
rect 6544 6384 6716 6434
rect 6480 6366 6544 6376
rect 6780 6384 7210 6434
rect 6716 6366 6780 6376
rect 5656 6304 5716 6314
rect 5158 6244 5656 6290
rect 5892 6304 5952 6314
rect 5716 6244 5892 6290
rect 6128 6304 6188 6314
rect 5952 6244 6128 6290
rect 6364 6304 6424 6314
rect 6188 6244 6364 6290
rect 6600 6304 6660 6314
rect 6424 6244 6600 6290
rect 6900 6292 6980 6302
rect 6900 6290 6910 6292
rect 6660 6244 6910 6290
rect 5158 6240 6910 6244
rect 3907 6234 6910 6240
rect 3907 6232 5532 6234
rect 6900 6232 6910 6234
rect 6970 6232 6980 6292
rect 3907 6231 3918 6232
rect 3836 6220 3918 6231
rect 4144 6230 4214 6232
rect 4380 6230 4450 6232
rect 4616 6230 4686 6232
rect 4852 6230 4922 6232
rect 5088 6230 5158 6232
rect 3615 6020 3893 6023
rect 4028 6020 4092 6024
rect 4264 6020 4328 6024
rect 4500 6020 4564 6024
rect 4736 6020 4800 6024
rect 4972 6020 5036 6024
rect 5208 6020 5272 6024
rect 3615 6014 5278 6020
rect 3615 5965 4028 6014
rect 3848 5962 4028 5965
rect 4092 5962 4264 6014
rect 4028 5944 4092 5954
rect 4328 5962 4500 6014
rect 4264 5944 4328 5954
rect 4564 5962 4736 6014
rect 4500 5944 4564 5954
rect 4800 5962 4972 6014
rect 4736 5944 4800 5954
rect 5036 5962 5208 6014
rect 4972 5944 5036 5954
rect 5272 5962 5278 6014
rect 5208 5944 5272 5954
rect 4144 5884 4214 5894
rect 3498 5876 3896 5878
rect 3491 5820 3500 5876
rect 3556 5824 4144 5876
rect 4380 5884 4450 5894
rect 4214 5824 4380 5876
rect 4616 5884 4686 5894
rect 4450 5824 4616 5876
rect 4852 5884 4922 5894
rect 4686 5824 4852 5876
rect 5088 5884 5158 5894
rect 4922 5824 5088 5876
rect 5375 5876 5446 6232
rect 6900 6222 6980 6232
rect 7155 6124 7210 6384
rect 5536 6022 5600 6024
rect 5772 6022 5836 6024
rect 6008 6022 6072 6024
rect 6244 6022 6308 6024
rect 6478 6022 6542 6024
rect 6716 6022 6780 6024
rect 7155 6022 7576 6124
rect 5524 6014 7576 6022
rect 7844 6114 7912 6122
rect 8360 6114 8428 6122
rect 8876 6114 8944 6122
rect 9392 6114 9460 6122
rect 9908 6114 9976 6122
rect 10424 6114 10492 6122
rect 10938 6114 11006 6122
rect 11456 6114 11524 6122
rect 11972 6114 12040 6122
rect 12488 6114 12556 6122
rect 13006 6114 13074 6122
rect 13242 6114 13318 6786
rect 13650 6114 13726 6786
rect 13984 6786 14430 6862
rect 13916 6766 13984 6776
rect 14498 6786 14948 6862
rect 14430 6766 14498 6776
rect 15016 6786 15464 6862
rect 14948 6766 15016 6776
rect 15532 6786 15980 6862
rect 15464 6766 15532 6776
rect 16048 6786 16498 6862
rect 15980 6766 16048 6776
rect 16566 6786 17010 6862
rect 16498 6766 16566 6776
rect 17078 6786 17528 6862
rect 17010 6766 17078 6776
rect 17596 6786 18042 6862
rect 17528 6766 17596 6776
rect 18110 6786 18560 6862
rect 18042 6766 18110 6776
rect 18628 6786 19076 6862
rect 18560 6766 18628 6776
rect 19144 6786 19160 6862
rect 19076 6766 19144 6776
rect 13916 6114 13984 6122
rect 14432 6114 14500 6124
rect 14948 6114 15016 6124
rect 15464 6114 15532 6124
rect 15980 6114 16048 6124
rect 16496 6114 16564 6124
rect 17012 6114 17080 6124
rect 17528 6114 17596 6124
rect 18044 6114 18112 6124
rect 18560 6114 18628 6124
rect 19076 6114 19144 6124
rect 7844 6112 14432 6114
rect 7912 6038 8360 6112
rect 7844 6016 7912 6026
rect 8428 6038 8876 6112
rect 8360 6016 8428 6026
rect 8944 6038 9392 6112
rect 8876 6016 8944 6026
rect 9460 6038 9908 6112
rect 9392 6016 9460 6026
rect 9976 6038 10424 6112
rect 9908 6016 9976 6026
rect 10492 6038 10938 6112
rect 10424 6016 10492 6026
rect 11006 6038 11456 6112
rect 10938 6016 11006 6026
rect 11524 6038 11972 6112
rect 11456 6016 11524 6026
rect 12040 6038 12488 6112
rect 11972 6016 12040 6026
rect 12556 6038 13006 6112
rect 12488 6016 12556 6026
rect 13074 6038 13916 6112
rect 13006 6016 13074 6026
rect 5524 5966 5536 6014
rect 5600 5966 5772 6014
rect 5536 5946 5600 5956
rect 5836 5966 6008 6014
rect 5772 5946 5836 5956
rect 6072 5966 6244 6014
rect 6008 5946 6072 5956
rect 6308 5966 6478 6014
rect 6244 5946 6308 5956
rect 6542 5966 6716 6014
rect 6478 5946 6542 5956
rect 6780 5967 7576 6014
rect 6780 5966 7002 5967
rect 7176 5964 7576 5967
rect 6716 5946 6780 5956
rect 5656 5886 5716 5896
rect 5158 5870 5534 5876
rect 5158 5826 5656 5870
rect 5892 5886 5952 5896
rect 5716 5826 5892 5870
rect 6128 5886 6188 5896
rect 5952 5826 6128 5870
rect 6366 5886 6426 5896
rect 6188 5826 6366 5870
rect 6600 5886 6660 5896
rect 6426 5826 6600 5870
rect 7278 5876 7335 5880
rect 6927 5871 7340 5876
rect 6927 5870 7278 5871
rect 6660 5826 7278 5870
rect 5158 5824 7278 5826
rect 3556 5820 7278 5824
rect 3498 5818 7278 5820
rect 4144 5814 4214 5818
rect 4380 5814 4450 5818
rect 4616 5814 4686 5818
rect 4852 5814 4922 5818
rect 5088 5814 5158 5818
rect 5272 5814 7278 5818
rect 7335 5814 7340 5871
rect 5375 5420 5446 5814
rect 6927 5809 7340 5814
rect 7278 5805 7335 5809
rect 5003 5257 5009 5420
rect 5172 5257 5650 5420
rect 5813 5257 5819 5420
rect 3873 4647 3879 4817
rect 4049 4647 4055 4817
rect 3879 4363 4049 4647
rect 469 4193 475 4363
rect 645 4195 4049 4363
rect 5311 4203 5505 5257
rect 7416 4392 7576 5964
rect 7844 5384 7912 5394
rect 8360 5384 8428 5394
rect 8878 5384 8946 5394
rect 9392 5384 9460 5394
rect 9908 5386 9976 5396
rect 7912 5308 8360 5384
rect 7844 5288 7912 5298
rect 8428 5308 8878 5384
rect 8360 5288 8428 5298
rect 8946 5308 9392 5384
rect 8878 5288 8946 5298
rect 9460 5308 9908 5384
rect 9392 5288 9460 5298
rect 10426 5386 10494 5396
rect 9976 5308 10426 5384
rect 9908 5290 9976 5300
rect 10940 5386 11008 5396
rect 10494 5308 10940 5384
rect 10426 5290 10494 5300
rect 11458 5386 11526 5396
rect 11008 5308 11458 5384
rect 10940 5290 11008 5300
rect 11972 5386 12040 5396
rect 11526 5308 11972 5384
rect 11458 5290 11526 5300
rect 12488 5386 12556 5396
rect 12040 5308 12488 5384
rect 11972 5290 12040 5300
rect 13006 5386 13074 5396
rect 12556 5308 13006 5384
rect 12488 5290 12556 5300
rect 13242 5384 13318 6038
rect 13650 5384 13726 6038
rect 13984 6038 14432 6112
rect 13916 6016 13984 6026
rect 14500 6038 14948 6114
rect 14432 6018 14500 6028
rect 15016 6038 15464 6114
rect 14948 6018 15016 6028
rect 15532 6038 15980 6114
rect 15464 6018 15532 6028
rect 16048 6038 16496 6114
rect 15980 6018 16048 6028
rect 16564 6038 17012 6114
rect 16496 6018 16564 6028
rect 17080 6038 17528 6114
rect 17012 6018 17080 6028
rect 17596 6038 18044 6114
rect 17528 6018 17596 6028
rect 18112 6038 18560 6114
rect 18044 6018 18112 6028
rect 18628 6038 19076 6114
rect 18560 6018 18628 6028
rect 19144 6038 19160 6114
rect 19076 6018 19144 6028
rect 13916 5386 13984 5396
rect 13074 5308 13916 5384
rect 13006 5290 13074 5300
rect 14434 5386 14502 5396
rect 13984 5308 14434 5384
rect 13916 5290 13984 5300
rect 14948 5386 15016 5396
rect 14502 5308 14948 5384
rect 14434 5290 14502 5300
rect 15464 5386 15532 5396
rect 15016 5308 15464 5384
rect 14948 5290 15016 5300
rect 15980 5386 16048 5396
rect 15532 5308 15980 5384
rect 15464 5290 15532 5300
rect 16496 5386 16564 5396
rect 16048 5308 16496 5384
rect 15980 5290 16048 5300
rect 17012 5386 17080 5396
rect 16564 5308 17012 5384
rect 16496 5290 16564 5300
rect 17528 5386 17596 5396
rect 17080 5308 17528 5384
rect 17012 5290 17080 5300
rect 18044 5386 18112 5396
rect 17596 5308 18044 5384
rect 17528 5290 17596 5300
rect 18560 5386 18628 5396
rect 18112 5308 18560 5384
rect 18044 5290 18112 5300
rect 19076 5386 19144 5396
rect 18628 5308 19076 5384
rect 18560 5290 18628 5300
rect 19144 5308 19160 5384
rect 19076 5290 19144 5300
rect 7416 4226 7576 4232
rect 645 4193 4036 4195
rect 5311 4009 6251 4203
rect 735 3853 1533 4002
rect 1682 3853 1688 4002
rect 746 2923 873 3853
rect 6057 3653 6251 4009
rect 8046 3790 8106 3800
rect 8282 3790 8342 3800
rect 8516 3790 8576 3800
rect 8752 3790 8812 3800
rect 8988 3790 9048 3800
rect 9224 3790 9284 3800
rect 9460 3790 9520 3800
rect 9696 3790 9756 3800
rect 9932 3790 9992 3800
rect 10168 3790 10228 3800
rect 8106 3714 8282 3790
rect 8046 3696 8106 3706
rect 8342 3714 8516 3790
rect 8282 3696 8342 3706
rect 8576 3714 8752 3790
rect 8516 3696 8576 3706
rect 8812 3714 8988 3790
rect 8752 3696 8812 3706
rect 9048 3714 9224 3790
rect 8988 3696 9048 3706
rect 9284 3714 9460 3790
rect 9224 3696 9284 3706
rect 9520 3714 9696 3790
rect 9460 3696 9520 3706
rect 9756 3714 9932 3790
rect 9696 3696 9756 3706
rect 9992 3714 10168 3790
rect 9932 3696 9992 3706
rect 10228 3714 10640 3790
rect 10168 3696 10228 3706
rect 1200 3522 1256 3532
rect 2116 3522 2172 3532
rect 3032 3522 3088 3532
rect 3948 3522 4004 3532
rect 4862 3522 4918 3528
rect 5778 3522 5834 3530
rect 6122 3522 6186 3653
rect 1182 3460 1200 3522
rect 1256 3460 2116 3522
rect 2172 3460 3032 3522
rect 3088 3460 3948 3522
rect 4004 3520 6200 3522
rect 4004 3518 5778 3520
rect 4004 3460 4862 3518
rect 1182 3458 4862 3460
rect 1200 3450 1256 3458
rect 2116 3450 2172 3458
rect 3032 3450 3088 3458
rect 3948 3450 4004 3458
rect 4918 3458 5778 3518
rect 5834 3458 6200 3520
rect 4862 3446 4918 3456
rect 5778 3448 5834 3458
rect 1652 3374 1722 3384
rect 2568 3374 2638 3384
rect 3482 3376 3552 3386
rect 1180 3318 1652 3374
rect 1722 3318 2568 3374
rect 2638 3320 3482 3374
rect 4400 3374 4470 3384
rect 5316 3374 5386 3384
rect 6998 3374 7004 3510
rect 7140 3480 7478 3510
rect 7922 3486 7990 3496
rect 7140 3404 7922 3480
rect 7140 3374 7478 3404
rect 8158 3486 8226 3496
rect 7990 3404 8158 3480
rect 7922 3392 7990 3402
rect 8396 3486 8464 3496
rect 8226 3404 8396 3480
rect 8158 3392 8226 3402
rect 8632 3486 8700 3496
rect 8464 3404 8632 3480
rect 8396 3392 8464 3402
rect 8868 3486 8936 3496
rect 8700 3404 8868 3480
rect 8632 3392 8700 3402
rect 9104 3486 9172 3496
rect 8936 3404 9104 3480
rect 8868 3392 8936 3402
rect 9340 3486 9408 3496
rect 9172 3404 9340 3480
rect 9104 3392 9172 3402
rect 9576 3488 9644 3498
rect 9408 3404 9576 3480
rect 9812 3488 9880 3498
rect 9644 3404 9812 3480
rect 10048 3488 10116 3498
rect 9880 3404 10048 3480
rect 10284 3488 10352 3498
rect 10116 3404 10284 3480
rect 9340 3392 9408 3402
rect 9576 3394 9644 3404
rect 9812 3394 9880 3404
rect 10048 3394 10116 3404
rect 10284 3394 10352 3404
rect 3552 3320 4400 3374
rect 2638 3318 4400 3320
rect 4470 3318 5316 3374
rect 5386 3318 6200 3374
rect 1180 3312 6200 3318
rect 1652 3308 1722 3312
rect 2568 3308 2638 3312
rect 3482 3310 3552 3312
rect 4400 3308 4470 3312
rect 5316 3308 5386 3312
rect 740 2796 746 2923
rect 873 2796 879 2923
rect 6137 2851 6199 3312
rect 6137 2783 6199 2789
rect 6348 2777 7003 2883
rect 7109 2777 7115 2883
rect 6348 2458 6454 2777
rect 7124 2458 7190 2460
rect 8042 2458 8108 2460
rect 8956 2458 9022 2460
rect 9872 2458 9938 2460
rect 10790 2458 10856 2460
rect 6348 2450 10856 2458
rect 6348 2404 7124 2450
rect 6348 2378 6454 2404
rect 7190 2404 8042 2450
rect 7124 2388 7190 2398
rect 8108 2404 8956 2450
rect 8042 2388 8108 2398
rect 9022 2404 9872 2450
rect 8956 2388 9022 2398
rect 9938 2404 10790 2450
rect 9872 2388 9938 2398
rect 10790 2388 10856 2398
rect 1190 2318 1260 2328
rect 912 2262 1190 2312
rect 2108 2320 2178 2330
rect 1260 2264 2108 2312
rect 3022 2320 3092 2330
rect 2178 2264 3022 2312
rect 3940 2320 4010 2330
rect 3092 2264 3940 2312
rect 4854 2320 4924 2330
rect 4010 2264 4854 2312
rect 5774 2320 5844 2330
rect 4924 2264 5774 2312
rect 6668 2314 6734 2324
rect 5844 2264 5860 2312
rect 1260 2262 5860 2264
rect 912 2252 5860 2262
rect 6660 2262 6668 2310
rect 7584 2314 7650 2324
rect 6734 2262 7584 2310
rect 8500 2314 8566 2324
rect 7650 2262 8500 2310
rect 9416 2314 9482 2324
rect 8566 2262 9416 2310
rect 10332 2314 10398 2324
rect 9482 2262 10332 2310
rect 11248 2314 11314 2324
rect 10398 2262 11248 2310
rect 11470 2310 11539 2318
rect 11314 2262 11542 2310
rect 6660 2256 11542 2262
rect 6668 2252 6734 2256
rect 7584 2252 7650 2256
rect 8500 2252 8566 2256
rect 9416 2252 9482 2256
rect 10332 2252 10398 2256
rect 11248 2252 11314 2256
rect 912 1480 972 2252
rect 11470 2051 11539 2256
rect 11470 1976 11539 1982
rect 1000 1494 1240 1504
rect 912 1420 1000 1480
rect 1000 1394 1240 1404
<< via2 >>
rect 3847 7487 3907 7547
rect 3847 7069 3907 7129
rect 6910 7482 6970 7542
rect 3847 6649 3907 6709
rect 6910 7064 6970 7124
rect 3847 6231 3907 6291
rect 6910 6652 6970 6712
rect 6910 6232 6970 6292
rect 3500 5820 3556 5876
rect 7278 5814 7335 5871
<< metal3 >>
rect 3842 7547 3912 7552
rect 3498 7487 3847 7547
rect 3907 7487 3912 7547
rect 3498 7129 3558 7487
rect 3842 7482 3912 7487
rect 6905 7542 6975 7547
rect 7273 7542 7340 7546
rect 6905 7482 6910 7542
rect 6970 7482 7340 7542
rect 6905 7477 6975 7482
rect 3842 7129 3912 7134
rect 3498 7069 3847 7129
rect 3907 7069 3912 7129
rect 3498 6709 3558 7069
rect 3842 7064 3912 7069
rect 6905 7124 6975 7129
rect 7273 7124 7340 7482
rect 6905 7064 6910 7124
rect 6970 7064 7340 7124
rect 6905 7059 6975 7064
rect 3842 6709 3912 6714
rect 3498 6649 3847 6709
rect 3907 6649 3912 6709
rect 3498 6291 3558 6649
rect 3842 6644 3912 6649
rect 6905 6712 6975 6717
rect 7273 6712 7340 7064
rect 6905 6652 6910 6712
rect 6970 6652 7340 6712
rect 6905 6647 6975 6652
rect 3842 6291 3912 6296
rect 3498 6231 3847 6291
rect 3907 6231 3912 6291
rect 3498 5881 3558 6231
rect 3842 6226 3912 6231
rect 6905 6292 6975 6297
rect 7273 6292 7340 6652
rect 6905 6232 6910 6292
rect 6970 6232 7340 6292
rect 6905 6227 6975 6232
rect 3495 5876 3561 5881
rect 3495 5820 3500 5876
rect 3556 5820 3561 5876
rect 3495 5815 3561 5820
rect 7273 5871 7340 6232
rect 7273 5814 7278 5871
rect 7335 5814 7340 5871
rect 7273 5809 7340 5814
use sky130_fd_pr__nfet_01v8_FMJ72H  XM1
timestamp 1713266475
transform 1 0 4651 0 1 6752
box -757 -1146 757 1146
use sky130_fd_pr__nfet_01v8_FMJ72H  XM2
timestamp 1713266475
transform 1 0 6159 0 1 6752
box -757 -1146 757 1146
use sky130_fd_pr__pfet_01v8_3H5TVM  XM3
timestamp 1713266475
transform 1 0 6410 0 1 9677
box -812 -319 812 319
use sky130_fd_pr__pfet_01v8_3H5TVM  XM4
timestamp 1713266475
transform 1 0 4454 0 1 9683
box -812 -319 812 319
use sky130_fd_pr__nfet_01v8_EPHDNF  XM5
timestamp 1713266475
transform 1 0 3517 0 1 3420
box -2457 -310 2457 310
use sky130_fd_pr__nfet_01v8_EPHDNF  XM6
timestamp 1713266475
transform 1 0 3517 0 1 2358
box -2457 -310 2457 310
use sky130_fd_pr__nfet_01v8_SMX62R  XM7
timestamp 1713266475
transform 1 0 9137 0 1 3602
box -1347 -410 1347 410
use sky130_fd_pr__nfet_01v8_EPHDNF  XM8
timestamp 1713266475
transform 1 0 8991 0 1 2356
box -2457 -310 2457 310
use sky130_fd_pr__pfet_01v8_P7N2DR  XM9
timestamp 1713266475
transform 1 0 10459 0 1 7343
box -2747 -2677 2747 2677
use sky130_fd_pr__pfet_01v8_P7N2DR  XM10
timestamp 1713266475
transform 1 0 16531 0 1 7343
box -2747 -2677 2747 2677
use sky130_fd_pr__nfet_01v8_EPHDNF  XM11
timestamp 1713266475
transform 1 0 14255 0 1 2358
box -2457 -310 2457 310
use sky130_fd_pr__nfet_01v8_V5FT3Q  XM12
timestamp 1713266475
transform 1 0 20546 0 1 3358
box -1312 -410 1312 410
use sky130_fd_pr__pfet_01v8_3HZ9VM  XM13
timestamp 1713266475
transform 1 0 20354 0 1 9245
box -296 -719 296 719
use sky130_fd_pr__nfet_01v8_EPHDNF  XM14
timestamp 1713266475
transform 1 0 19417 0 1 2358
box -2457 -310 2457 310
use sky130_fd_pr__nfet_01v8_GSBCLJ  XM15
timestamp 1713266475
transform 1 0 21111 0 1 5197
box -647 -1119 647 1119
use sky130_fd_pr__pfet_01v8_3HZ9VM  XM16
timestamp 1713266475
transform 1 0 21446 0 1 9243
box -296 -719 296 719
use sky130_fd_pr__pfet_01v8_BDVWJN  XM17
timestamp 1713266475
transform 1 0 21123 0 1 7365
box -647 -719 647 719
use sky130_fd_pr__res_xhigh_po_0p35_RF5GSL  XR1
timestamp 1713266475
transform 1 0 1553 0 1 6300
box -201 -1382 201 1382
use sky130_fd_pr__res_xhigh_po_0p35_RF5GSL  XR2
timestamp 1713266475
transform 1 0 1161 0 1 6300
box -201 -1382 201 1382
use sky130_fd_pr__res_xhigh_po_0p35_RF5GSL  XR3
timestamp 1713266475
transform 1 0 1947 0 1 6300
box -201 -1382 201 1382
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR4
timestamp 1713266475
transform 1 0 2345 0 1 6500
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR5
timestamp 1713266475
transform 1 0 3143 0 1 6500
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR6
timestamp 1713266475
transform 1 0 2749 0 1 6500
box -201 -1582 201 1582
<< labels >>
flabel metal1 106 1246 306 1446 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 22378 6402 22578 6602 0 FreeSans 256 0 0 0 z
port 2 nsew
flabel metal1 22380 4698 22580 4898 0 FreeSans 256 0 0 0 x
port 5 nsew
flabel metal1 98 4186 298 4386 0 FreeSans 256 0 0 0 y
port 3 nsew
flabel metal1 102 8284 302 8484 0 FreeSans 256 0 0 0 ref
port 4 nsew
flabel metal1 92 10506 292 10706 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 3428 3864 6574 4072 0 FreeSans 1600 0 0 0 G2
flabel metal1 5370 9488 5476 9876 0 FreeSans 1600 0 0 0 G1
flabel metal2 7057 7638 7203 8921 0 FreeSans 1600 0 0 0 D1
flabel metal2 5172 5257 5650 5420 0 FreeSans 1600 0 0 0 B1
<< end >>
