magic
tech sky130A
magscale 1 2
timestamp 1713266475
<< pwell >>
rect -2457 -310 2457 310
<< nmos >>
rect -2261 -100 -1861 100
rect -1803 -100 -1403 100
rect -1345 -100 -945 100
rect -887 -100 -487 100
rect -429 -100 -29 100
rect 29 -100 429 100
rect 487 -100 887 100
rect 945 -100 1345 100
rect 1403 -100 1803 100
rect 1861 -100 2261 100
<< ndiff >>
rect -2319 88 -2261 100
rect -2319 -88 -2307 88
rect -2273 -88 -2261 88
rect -2319 -100 -2261 -88
rect -1861 88 -1803 100
rect -1861 -88 -1849 88
rect -1815 -88 -1803 88
rect -1861 -100 -1803 -88
rect -1403 88 -1345 100
rect -1403 -88 -1391 88
rect -1357 -88 -1345 88
rect -1403 -100 -1345 -88
rect -945 88 -887 100
rect -945 -88 -933 88
rect -899 -88 -887 88
rect -945 -100 -887 -88
rect -487 88 -429 100
rect -487 -88 -475 88
rect -441 -88 -429 88
rect -487 -100 -429 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 429 88 487 100
rect 429 -88 441 88
rect 475 -88 487 88
rect 429 -100 487 -88
rect 887 88 945 100
rect 887 -88 899 88
rect 933 -88 945 88
rect 887 -100 945 -88
rect 1345 88 1403 100
rect 1345 -88 1357 88
rect 1391 -88 1403 88
rect 1345 -100 1403 -88
rect 1803 88 1861 100
rect 1803 -88 1815 88
rect 1849 -88 1861 88
rect 1803 -100 1861 -88
rect 2261 88 2319 100
rect 2261 -88 2273 88
rect 2307 -88 2319 88
rect 2261 -100 2319 -88
<< ndiffc >>
rect -2307 -88 -2273 88
rect -1849 -88 -1815 88
rect -1391 -88 -1357 88
rect -933 -88 -899 88
rect -475 -88 -441 88
rect -17 -88 17 88
rect 441 -88 475 88
rect 899 -88 933 88
rect 1357 -88 1391 88
rect 1815 -88 1849 88
rect 2273 -88 2307 88
<< psubdiff >>
rect -2421 240 -2325 274
rect 2325 240 2421 274
rect -2421 178 -2387 240
rect 2387 178 2421 240
rect -2421 -240 -2387 -178
rect 2387 -240 2421 -178
rect -2421 -274 -2325 -240
rect 2325 -274 2421 -240
<< psubdiffcont >>
rect -2325 240 2325 274
rect -2421 -178 -2387 178
rect 2387 -178 2421 178
rect -2325 -274 2325 -240
<< poly >>
rect -2261 172 -1861 188
rect -2261 138 -2245 172
rect -1877 138 -1861 172
rect -2261 100 -1861 138
rect -1803 172 -1403 188
rect -1803 138 -1787 172
rect -1419 138 -1403 172
rect -1803 100 -1403 138
rect -1345 172 -945 188
rect -1345 138 -1329 172
rect -961 138 -945 172
rect -1345 100 -945 138
rect -887 172 -487 188
rect -887 138 -871 172
rect -503 138 -487 172
rect -887 100 -487 138
rect -429 172 -29 188
rect -429 138 -413 172
rect -45 138 -29 172
rect -429 100 -29 138
rect 29 172 429 188
rect 29 138 45 172
rect 413 138 429 172
rect 29 100 429 138
rect 487 172 887 188
rect 487 138 503 172
rect 871 138 887 172
rect 487 100 887 138
rect 945 172 1345 188
rect 945 138 961 172
rect 1329 138 1345 172
rect 945 100 1345 138
rect 1403 172 1803 188
rect 1403 138 1419 172
rect 1787 138 1803 172
rect 1403 100 1803 138
rect 1861 172 2261 188
rect 1861 138 1877 172
rect 2245 138 2261 172
rect 1861 100 2261 138
rect -2261 -138 -1861 -100
rect -2261 -172 -2245 -138
rect -1877 -172 -1861 -138
rect -2261 -188 -1861 -172
rect -1803 -138 -1403 -100
rect -1803 -172 -1787 -138
rect -1419 -172 -1403 -138
rect -1803 -188 -1403 -172
rect -1345 -138 -945 -100
rect -1345 -172 -1329 -138
rect -961 -172 -945 -138
rect -1345 -188 -945 -172
rect -887 -138 -487 -100
rect -887 -172 -871 -138
rect -503 -172 -487 -138
rect -887 -188 -487 -172
rect -429 -138 -29 -100
rect -429 -172 -413 -138
rect -45 -172 -29 -138
rect -429 -188 -29 -172
rect 29 -138 429 -100
rect 29 -172 45 -138
rect 413 -172 429 -138
rect 29 -188 429 -172
rect 487 -138 887 -100
rect 487 -172 503 -138
rect 871 -172 887 -138
rect 487 -188 887 -172
rect 945 -138 1345 -100
rect 945 -172 961 -138
rect 1329 -172 1345 -138
rect 945 -188 1345 -172
rect 1403 -138 1803 -100
rect 1403 -172 1419 -138
rect 1787 -172 1803 -138
rect 1403 -188 1803 -172
rect 1861 -138 2261 -100
rect 1861 -172 1877 -138
rect 2245 -172 2261 -138
rect 1861 -188 2261 -172
<< polycont >>
rect -2245 138 -1877 172
rect -1787 138 -1419 172
rect -1329 138 -961 172
rect -871 138 -503 172
rect -413 138 -45 172
rect 45 138 413 172
rect 503 138 871 172
rect 961 138 1329 172
rect 1419 138 1787 172
rect 1877 138 2245 172
rect -2245 -172 -1877 -138
rect -1787 -172 -1419 -138
rect -1329 -172 -961 -138
rect -871 -172 -503 -138
rect -413 -172 -45 -138
rect 45 -172 413 -138
rect 503 -172 871 -138
rect 961 -172 1329 -138
rect 1419 -172 1787 -138
rect 1877 -172 2245 -138
<< locali >>
rect -2421 240 -2325 274
rect 2325 240 2421 274
rect -2421 178 -2387 240
rect 2387 178 2421 240
rect -2261 138 -2245 172
rect -1877 138 -1861 172
rect -1803 138 -1787 172
rect -1419 138 -1403 172
rect -1345 138 -1329 172
rect -961 138 -945 172
rect -887 138 -871 172
rect -503 138 -487 172
rect -429 138 -413 172
rect -45 138 -29 172
rect 29 138 45 172
rect 413 138 429 172
rect 487 138 503 172
rect 871 138 887 172
rect 945 138 961 172
rect 1329 138 1345 172
rect 1403 138 1419 172
rect 1787 138 1803 172
rect 1861 138 1877 172
rect 2245 138 2261 172
rect -2307 88 -2273 104
rect -2307 -104 -2273 -88
rect -1849 88 -1815 104
rect -1849 -104 -1815 -88
rect -1391 88 -1357 104
rect -1391 -104 -1357 -88
rect -933 88 -899 104
rect -933 -104 -899 -88
rect -475 88 -441 104
rect -475 -104 -441 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 441 88 475 104
rect 441 -104 475 -88
rect 899 88 933 104
rect 899 -104 933 -88
rect 1357 88 1391 104
rect 1357 -104 1391 -88
rect 1815 88 1849 104
rect 1815 -104 1849 -88
rect 2273 88 2307 104
rect 2273 -104 2307 -88
rect -2261 -172 -2245 -138
rect -1877 -172 -1861 -138
rect -1803 -172 -1787 -138
rect -1419 -172 -1403 -138
rect -1345 -172 -1329 -138
rect -961 -172 -945 -138
rect -887 -172 -871 -138
rect -503 -172 -487 -138
rect -429 -172 -413 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 413 -172 429 -138
rect 487 -172 503 -138
rect 871 -172 887 -138
rect 945 -172 961 -138
rect 1329 -172 1345 -138
rect 1403 -172 1419 -138
rect 1787 -172 1803 -138
rect 1861 -172 1877 -138
rect 2245 -172 2261 -138
rect -2421 -240 -2387 -178
rect 2387 -240 2421 -178
rect -2421 -274 -2325 -240
rect 2325 -274 2421 -240
<< viali >>
rect -2245 138 -1877 172
rect -1787 138 -1419 172
rect -1329 138 -961 172
rect -871 138 -503 172
rect -413 138 -45 172
rect 45 138 413 172
rect 503 138 871 172
rect 961 138 1329 172
rect 1419 138 1787 172
rect 1877 138 2245 172
rect -2307 -88 -2273 88
rect -1849 -88 -1815 88
rect -1391 -88 -1357 88
rect -933 -88 -899 88
rect -475 -88 -441 88
rect -17 -88 17 88
rect 441 -88 475 88
rect 899 -88 933 88
rect 1357 -88 1391 88
rect 1815 -88 1849 88
rect 2273 -88 2307 88
rect -2245 -172 -1877 -138
rect -1787 -172 -1419 -138
rect -1329 -172 -961 -138
rect -871 -172 -503 -138
rect -413 -172 -45 -138
rect 45 -172 413 -138
rect 503 -172 871 -138
rect 961 -172 1329 -138
rect 1419 -172 1787 -138
rect 1877 -172 2245 -138
<< metal1 >>
rect -2257 172 -1865 178
rect -2257 138 -2245 172
rect -1877 138 -1865 172
rect -2257 132 -1865 138
rect -1799 172 -1407 178
rect -1799 138 -1787 172
rect -1419 138 -1407 172
rect -1799 132 -1407 138
rect -1341 172 -949 178
rect -1341 138 -1329 172
rect -961 138 -949 172
rect -1341 132 -949 138
rect -883 172 -491 178
rect -883 138 -871 172
rect -503 138 -491 172
rect -883 132 -491 138
rect -425 172 -33 178
rect -425 138 -413 172
rect -45 138 -33 172
rect -425 132 -33 138
rect 33 172 425 178
rect 33 138 45 172
rect 413 138 425 172
rect 33 132 425 138
rect 491 172 883 178
rect 491 138 503 172
rect 871 138 883 172
rect 491 132 883 138
rect 949 172 1341 178
rect 949 138 961 172
rect 1329 138 1341 172
rect 949 132 1341 138
rect 1407 172 1799 178
rect 1407 138 1419 172
rect 1787 138 1799 172
rect 1407 132 1799 138
rect 1865 172 2257 178
rect 1865 138 1877 172
rect 2245 138 2257 172
rect 1865 132 2257 138
rect -2313 88 -2267 100
rect -2313 -88 -2307 88
rect -2273 -88 -2267 88
rect -2313 -100 -2267 -88
rect -1855 88 -1809 100
rect -1855 -88 -1849 88
rect -1815 -88 -1809 88
rect -1855 -100 -1809 -88
rect -1397 88 -1351 100
rect -1397 -88 -1391 88
rect -1357 -88 -1351 88
rect -1397 -100 -1351 -88
rect -939 88 -893 100
rect -939 -88 -933 88
rect -899 -88 -893 88
rect -939 -100 -893 -88
rect -481 88 -435 100
rect -481 -88 -475 88
rect -441 -88 -435 88
rect -481 -100 -435 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 435 88 481 100
rect 435 -88 441 88
rect 475 -88 481 88
rect 435 -100 481 -88
rect 893 88 939 100
rect 893 -88 899 88
rect 933 -88 939 88
rect 893 -100 939 -88
rect 1351 88 1397 100
rect 1351 -88 1357 88
rect 1391 -88 1397 88
rect 1351 -100 1397 -88
rect 1809 88 1855 100
rect 1809 -88 1815 88
rect 1849 -88 1855 88
rect 1809 -100 1855 -88
rect 2267 88 2313 100
rect 2267 -88 2273 88
rect 2307 -88 2313 88
rect 2267 -100 2313 -88
rect -2257 -138 -1865 -132
rect -2257 -172 -2245 -138
rect -1877 -172 -1865 -138
rect -2257 -178 -1865 -172
rect -1799 -138 -1407 -132
rect -1799 -172 -1787 -138
rect -1419 -172 -1407 -138
rect -1799 -178 -1407 -172
rect -1341 -138 -949 -132
rect -1341 -172 -1329 -138
rect -961 -172 -949 -138
rect -1341 -178 -949 -172
rect -883 -138 -491 -132
rect -883 -172 -871 -138
rect -503 -172 -491 -138
rect -883 -178 -491 -172
rect -425 -138 -33 -132
rect -425 -172 -413 -138
rect -45 -172 -33 -138
rect -425 -178 -33 -172
rect 33 -138 425 -132
rect 33 -172 45 -138
rect 413 -172 425 -138
rect 33 -178 425 -172
rect 491 -138 883 -132
rect 491 -172 503 -138
rect 871 -172 883 -138
rect 491 -178 883 -172
rect 949 -138 1341 -132
rect 949 -172 961 -138
rect 1329 -172 1341 -138
rect 949 -178 1341 -172
rect 1407 -138 1799 -132
rect 1407 -172 1419 -138
rect 1787 -172 1799 -138
rect 1407 -178 1799 -172
rect 1865 -138 2257 -132
rect 1865 -172 1877 -138
rect 2245 -172 2257 -138
rect 1865 -178 2257 -172
<< properties >>
string FIXED_BBOX -2404 -257 2404 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 2.0 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
