magic
tech sky130A
magscale 1 2
timestamp 1713521240
<< metal1 >>
rect 20546 32466 21015 32551
rect 20546 32166 20630 32466
rect 20930 32166 21015 32466
rect 20546 29064 21015 32166
rect 29800 32522 30240 32592
rect 29800 32222 29870 32522
rect 30170 32222 30240 32522
rect 23627 29561 23633 29739
rect 23811 29561 23817 29739
rect 27745 29720 27918 29721
rect 23633 29111 23811 29561
rect 27740 29549 27746 29720
rect 27917 29549 27923 29720
rect 27745 29122 27918 29549
rect 29800 28912 30240 32222
rect 24672 6508 24833 7052
rect 24666 6347 24672 6508
rect 24833 6347 24839 6508
rect 25824 6414 26008 7046
rect 25824 6265 25842 6414
rect 25991 6265 26008 6414
rect 25824 6247 26008 6265
<< via1 >>
rect 20630 32166 20930 32466
rect 29870 32222 30170 32522
rect 23633 29561 23811 29739
rect 27746 29549 27917 29720
rect 24672 6347 24833 6508
rect 25842 6265 25991 6414
<< metal2 >>
rect 29870 33727 30170 33732
rect 29866 33437 29875 33727
rect 30165 33437 30174 33727
rect 20630 33009 20930 33014
rect 20626 32719 20635 33009
rect 20925 32719 20934 33009
rect 20630 32466 20930 32719
rect 29870 32522 30170 33437
rect 29870 32216 30170 32222
rect 20630 32160 20930 32166
rect 23633 29982 23811 29987
rect 23629 29814 23638 29982
rect 23806 29814 23815 29982
rect 27746 29971 27917 29976
rect 23633 29739 23811 29814
rect 27742 29810 27751 29971
rect 27912 29810 27921 29971
rect 23633 29555 23811 29561
rect 27746 29720 27917 29810
rect 27746 29543 27917 29549
rect 24672 6508 24833 6514
rect 24672 6187 24833 6347
rect 25842 6414 25991 6420
rect 25842 6197 25991 6265
rect 24668 6036 24677 6187
rect 24828 6036 24837 6187
rect 25838 6058 25847 6197
rect 25986 6058 25995 6197
rect 25842 6053 25991 6058
rect 24672 6031 24833 6036
<< via2 >>
rect 29875 33437 30165 33727
rect 20635 32719 20925 33009
rect 23638 29814 23806 29982
rect 27751 29810 27912 29971
rect 24677 6036 24828 6187
rect 25847 6058 25986 6197
<< metal3 >>
rect 6595 35462 6893 35467
rect 6594 35461 30170 35462
rect 6594 35163 6595 35461
rect 6893 35163 30170 35461
rect 6594 35162 30170 35163
rect 6595 35157 6893 35162
rect 20630 33737 20930 33738
rect 20625 33439 20631 33737
rect 20929 33439 20935 33737
rect 29870 33727 30170 35162
rect 20630 33009 20930 33439
rect 29870 33437 29875 33727
rect 30165 33437 30170 33727
rect 29870 33432 30170 33437
rect 20630 32719 20635 33009
rect 20925 32719 20930 33009
rect 20630 32714 20930 32719
rect 27746 30241 27917 30242
rect 23633 30234 23811 30235
rect 23628 30058 23634 30234
rect 23810 30058 23816 30234
rect 27741 30072 27747 30241
rect 27916 30072 27922 30241
rect 23633 29982 23811 30058
rect 23633 29814 23638 29982
rect 23806 29814 23811 29982
rect 23633 29809 23811 29814
rect 27746 29971 27917 30072
rect 27746 29810 27751 29971
rect 27912 29810 27917 29971
rect 27746 29805 27917 29810
rect 25842 6197 25991 6202
rect 24672 6187 24833 6192
rect 24672 6036 24677 6187
rect 24828 6036 24833 6187
rect 24672 5831 24833 6036
rect 25842 6058 25847 6197
rect 25986 6058 25991 6197
rect 25842 5858 25991 6058
rect 24672 5672 24673 5831
rect 24832 5672 24833 5831
rect 25837 5711 25843 5858
rect 25990 5711 25996 5858
rect 25842 5710 25991 5711
rect 24672 5671 24833 5672
rect 24673 5666 24832 5671
<< via3 >>
rect 6595 35163 6893 35461
rect 20631 33439 20929 33737
rect 23634 30058 23810 30234
rect 27747 30072 27916 30241
rect 24673 5672 24832 5831
rect 25843 5711 25990 5858
<< metal4 >>
rect 798 44750 858 45152
rect 1534 44750 1594 45152
rect 2270 44750 2330 45152
rect 3006 44750 3066 45152
rect 3742 44750 3802 45152
rect 4478 44750 4538 45152
rect 5214 44750 5274 45152
rect 5950 44750 6010 45152
rect 6686 44750 6746 45152
rect 7422 44750 7482 45152
rect 8158 44750 8218 45152
rect 8894 44750 8954 45152
rect 9630 44750 9690 45152
rect 10366 44750 10426 45152
rect 11102 44750 11162 45152
rect 11838 44750 11898 45152
rect 12574 44750 12634 45152
rect 13310 44750 13370 45152
rect 14046 44750 14106 45152
rect 14782 44750 14842 45152
rect 15518 44750 15578 45152
rect 16254 44750 16314 45152
rect 16990 44750 17050 45152
rect 17726 44750 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 762 44418 17786 44750
rect 200 35462 500 44152
rect 200 35461 6894 35462
rect 200 35163 6595 35461
rect 6893 35163 6894 35461
rect 200 35162 6894 35163
rect 200 1000 500 35162
rect 9800 33738 10100 44418
rect 17726 44416 17786 44418
rect 9800 33737 20930 33738
rect 9800 33439 20631 33737
rect 20929 33439 20930 33737
rect 9800 33438 20930 33439
rect 9800 1000 10100 33438
rect 16618 31293 27917 31464
rect 16618 4238 16789 31293
rect 18035 30355 23811 30533
rect 18064 5125 18184 30355
rect 23633 30234 23811 30355
rect 23633 30058 23634 30234
rect 23810 30058 23811 30234
rect 27746 30241 27917 31293
rect 27746 30072 27747 30241
rect 27916 30072 27917 30241
rect 27746 30071 27917 30072
rect 23633 30057 23811 30058
rect 25842 5858 31447 5859
rect 24672 5831 24833 5832
rect 24672 5672 24673 5831
rect 24832 5672 24833 5831
rect 25842 5711 25843 5858
rect 25990 5711 31447 5858
rect 25842 5710 31447 5711
rect 18064 5003 22601 5125
rect 18064 5000 18184 5003
rect 16618 4118 18184 4238
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 202
rect 18064 0 18184 4118
rect 22479 2648 22601 5003
rect 24672 4843 24833 5672
rect 24672 4682 27037 4843
rect 22479 -1 22602 2648
rect 26896 0 27016 4682
rect 31312 0 31432 5710
use VCII-final  VCII-final_0
timestamp 1713478763
transform 0 1 19454 -1 0 29407
box 10 1078 22641 10794
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
