magic
tech sky130A
magscale 1 2
timestamp 1713335455
<< error_s >>
rect 20758 7946 20816 7952
rect 20950 7946 21008 7952
rect 21142 7946 21200 7952
rect 21334 7946 21392 7952
rect 21526 7946 21584 7952
rect 20758 7912 20770 7946
rect 20950 7912 20962 7946
rect 21142 7912 21154 7946
rect 21334 7912 21346 7946
rect 21526 7912 21538 7946
rect 20758 7906 20816 7912
rect 20950 7906 21008 7912
rect 21142 7906 21200 7912
rect 21334 7906 21392 7912
rect 21526 7906 21584 7912
rect 4091 7760 4149 7766
rect 4209 7760 4267 7766
rect 4327 7760 4385 7766
rect 4445 7760 4503 7766
rect 4563 7760 4621 7766
rect 4681 7760 4739 7766
rect 4799 7760 4857 7766
rect 4917 7760 4975 7766
rect 5035 7760 5093 7766
rect 5153 7760 5211 7766
rect 5599 7760 5657 7766
rect 5717 7760 5775 7766
rect 5835 7760 5893 7766
rect 5953 7760 6011 7766
rect 6071 7760 6129 7766
rect 6189 7760 6247 7766
rect 6307 7760 6365 7766
rect 6425 7760 6483 7766
rect 6543 7760 6601 7766
rect 6661 7760 6719 7766
rect 4091 7726 4103 7760
rect 4209 7726 4221 7760
rect 4327 7726 4339 7760
rect 4445 7726 4457 7760
rect 4563 7726 4575 7760
rect 4681 7726 4693 7760
rect 4799 7726 4811 7760
rect 4917 7726 4929 7760
rect 5035 7726 5047 7760
rect 5153 7726 5165 7760
rect 5599 7726 5611 7760
rect 5717 7726 5729 7760
rect 5835 7726 5847 7760
rect 5953 7726 5965 7760
rect 6071 7726 6083 7760
rect 6189 7726 6201 7760
rect 6307 7726 6319 7760
rect 6425 7726 6437 7760
rect 6543 7726 6555 7760
rect 6661 7726 6673 7760
rect 4091 7720 4149 7726
rect 4209 7720 4267 7726
rect 4327 7720 4385 7726
rect 4445 7720 4503 7726
rect 4563 7720 4621 7726
rect 4681 7720 4739 7726
rect 4799 7720 4857 7726
rect 4917 7720 4975 7726
rect 5035 7720 5093 7726
rect 5153 7720 5211 7726
rect 5599 7720 5657 7726
rect 5717 7720 5775 7726
rect 5835 7720 5893 7726
rect 5953 7720 6011 7726
rect 6071 7720 6129 7726
rect 6189 7720 6247 7726
rect 6307 7720 6365 7726
rect 6425 7720 6483 7726
rect 6543 7720 6601 7726
rect 6661 7720 6719 7726
rect 4091 7450 4149 7456
rect 4209 7450 4267 7456
rect 4327 7450 4385 7456
rect 4445 7450 4503 7456
rect 4563 7450 4621 7456
rect 4681 7450 4739 7456
rect 4799 7450 4857 7456
rect 4917 7450 4975 7456
rect 5035 7450 5093 7456
rect 5153 7450 5211 7456
rect 5599 7450 5657 7456
rect 5717 7450 5775 7456
rect 5835 7450 5893 7456
rect 5953 7450 6011 7456
rect 6071 7450 6129 7456
rect 6189 7450 6247 7456
rect 6307 7450 6365 7456
rect 6425 7450 6483 7456
rect 6543 7450 6601 7456
rect 6661 7450 6719 7456
rect 4091 7416 4103 7450
rect 4209 7416 4221 7450
rect 4327 7416 4339 7450
rect 4445 7416 4457 7450
rect 4563 7416 4575 7450
rect 4681 7416 4693 7450
rect 4799 7416 4811 7450
rect 4917 7416 4929 7450
rect 5035 7416 5047 7450
rect 5153 7416 5165 7450
rect 5599 7416 5611 7450
rect 5717 7416 5729 7450
rect 5835 7416 5847 7450
rect 5953 7416 5965 7450
rect 6071 7416 6083 7450
rect 6189 7416 6201 7450
rect 6307 7416 6319 7450
rect 6425 7416 6437 7450
rect 6543 7416 6555 7450
rect 6661 7416 6673 7450
rect 4091 7410 4149 7416
rect 4209 7410 4267 7416
rect 4327 7410 4385 7416
rect 4445 7410 4503 7416
rect 4563 7410 4621 7416
rect 4681 7410 4739 7416
rect 4799 7410 4857 7416
rect 4917 7410 4975 7416
rect 5035 7410 5093 7416
rect 5153 7410 5211 7416
rect 5599 7410 5657 7416
rect 5717 7410 5775 7416
rect 5835 7410 5893 7416
rect 5953 7410 6011 7416
rect 6071 7410 6129 7416
rect 6189 7410 6247 7416
rect 6307 7410 6365 7416
rect 6425 7410 6483 7416
rect 6543 7410 6601 7416
rect 6661 7410 6719 7416
rect 4091 7342 4149 7348
rect 4209 7342 4267 7348
rect 4327 7342 4385 7348
rect 4445 7342 4503 7348
rect 4563 7342 4621 7348
rect 4681 7342 4739 7348
rect 4799 7342 4857 7348
rect 4917 7342 4975 7348
rect 5035 7342 5093 7348
rect 5153 7342 5211 7348
rect 5599 7342 5657 7348
rect 5717 7342 5775 7348
rect 5835 7342 5893 7348
rect 5953 7342 6011 7348
rect 6071 7342 6129 7348
rect 6189 7342 6247 7348
rect 6307 7342 6365 7348
rect 6425 7342 6483 7348
rect 6543 7342 6601 7348
rect 6661 7342 6719 7348
rect 4091 7308 4103 7342
rect 4209 7308 4221 7342
rect 4327 7308 4339 7342
rect 4445 7308 4457 7342
rect 4563 7308 4575 7342
rect 4681 7308 4693 7342
rect 4799 7308 4811 7342
rect 4917 7308 4929 7342
rect 5035 7308 5047 7342
rect 5153 7308 5165 7342
rect 5599 7308 5611 7342
rect 5717 7308 5729 7342
rect 5835 7308 5847 7342
rect 5953 7308 5965 7342
rect 6071 7308 6083 7342
rect 6189 7308 6201 7342
rect 6307 7308 6319 7342
rect 6425 7308 6437 7342
rect 6543 7308 6555 7342
rect 6661 7308 6673 7342
rect 4091 7302 4149 7308
rect 4209 7302 4267 7308
rect 4327 7302 4385 7308
rect 4445 7302 4503 7308
rect 4563 7302 4621 7308
rect 4681 7302 4739 7308
rect 4799 7302 4857 7308
rect 4917 7302 4975 7308
rect 5035 7302 5093 7308
rect 5153 7302 5211 7308
rect 5599 7302 5657 7308
rect 5717 7302 5775 7308
rect 5835 7302 5893 7308
rect 5953 7302 6011 7308
rect 6071 7302 6129 7308
rect 6189 7302 6247 7308
rect 6307 7302 6365 7308
rect 6425 7302 6483 7308
rect 6543 7302 6601 7308
rect 6661 7302 6719 7308
rect 4091 7032 4149 7038
rect 4209 7032 4267 7038
rect 4327 7032 4385 7038
rect 4445 7032 4503 7038
rect 4563 7032 4621 7038
rect 4681 7032 4739 7038
rect 4799 7032 4857 7038
rect 4917 7032 4975 7038
rect 5035 7032 5093 7038
rect 5153 7032 5211 7038
rect 5599 7032 5657 7038
rect 5717 7032 5775 7038
rect 5835 7032 5893 7038
rect 5953 7032 6011 7038
rect 6071 7032 6129 7038
rect 6189 7032 6247 7038
rect 6307 7032 6365 7038
rect 6425 7032 6483 7038
rect 6543 7032 6601 7038
rect 6661 7032 6719 7038
rect 4091 6998 4103 7032
rect 4209 6998 4221 7032
rect 4327 6998 4339 7032
rect 4445 6998 4457 7032
rect 4563 6998 4575 7032
rect 4681 6998 4693 7032
rect 4799 6998 4811 7032
rect 4917 6998 4929 7032
rect 5035 6998 5047 7032
rect 5153 6998 5165 7032
rect 5599 6998 5611 7032
rect 5717 6998 5729 7032
rect 5835 6998 5847 7032
rect 5953 6998 5965 7032
rect 6071 6998 6083 7032
rect 6189 6998 6201 7032
rect 6307 6998 6319 7032
rect 6425 6998 6437 7032
rect 6543 6998 6555 7032
rect 6661 6998 6673 7032
rect 4091 6992 4149 6998
rect 4209 6992 4267 6998
rect 4327 6992 4385 6998
rect 4445 6992 4503 6998
rect 4563 6992 4621 6998
rect 4681 6992 4739 6998
rect 4799 6992 4857 6998
rect 4917 6992 4975 6998
rect 5035 6992 5093 6998
rect 5153 6992 5211 6998
rect 5599 6992 5657 6998
rect 5717 6992 5775 6998
rect 5835 6992 5893 6998
rect 5953 6992 6011 6998
rect 6071 6992 6129 6998
rect 6189 6992 6247 6998
rect 6307 6992 6365 6998
rect 6425 6992 6483 6998
rect 6543 6992 6601 6998
rect 6661 6992 6719 6998
rect 4091 6924 4149 6930
rect 4209 6924 4267 6930
rect 4327 6924 4385 6930
rect 4445 6924 4503 6930
rect 4563 6924 4621 6930
rect 4681 6924 4739 6930
rect 4799 6924 4857 6930
rect 4917 6924 4975 6930
rect 5035 6924 5093 6930
rect 5153 6924 5211 6930
rect 5599 6924 5657 6930
rect 5717 6924 5775 6930
rect 5835 6924 5893 6930
rect 5953 6924 6011 6930
rect 6071 6924 6129 6930
rect 6189 6924 6247 6930
rect 6307 6924 6365 6930
rect 6425 6924 6483 6930
rect 6543 6924 6601 6930
rect 6661 6924 6719 6930
rect 4091 6890 4103 6924
rect 4209 6890 4221 6924
rect 4327 6890 4339 6924
rect 4445 6890 4457 6924
rect 4563 6890 4575 6924
rect 4681 6890 4693 6924
rect 4799 6890 4811 6924
rect 4917 6890 4929 6924
rect 5035 6890 5047 6924
rect 5153 6890 5165 6924
rect 5599 6890 5611 6924
rect 5717 6890 5729 6924
rect 5835 6890 5847 6924
rect 5953 6890 5965 6924
rect 6071 6890 6083 6924
rect 6189 6890 6201 6924
rect 6307 6890 6319 6924
rect 6425 6890 6437 6924
rect 6543 6890 6555 6924
rect 6661 6890 6673 6924
rect 4091 6884 4149 6890
rect 4209 6884 4267 6890
rect 4327 6884 4385 6890
rect 4445 6884 4503 6890
rect 4563 6884 4621 6890
rect 4681 6884 4739 6890
rect 4799 6884 4857 6890
rect 4917 6884 4975 6890
rect 5035 6884 5093 6890
rect 5153 6884 5211 6890
rect 5599 6884 5657 6890
rect 5717 6884 5775 6890
rect 5835 6884 5893 6890
rect 5953 6884 6011 6890
rect 6071 6884 6129 6890
rect 6189 6884 6247 6890
rect 6307 6884 6365 6890
rect 6425 6884 6483 6890
rect 6543 6884 6601 6890
rect 6661 6884 6719 6890
rect 20662 6818 20720 6824
rect 20854 6818 20912 6824
rect 21046 6818 21104 6824
rect 21238 6818 21296 6824
rect 21430 6818 21488 6824
rect 20662 6784 20674 6818
rect 20854 6784 20866 6818
rect 21046 6784 21058 6818
rect 21238 6784 21250 6818
rect 21430 6784 21442 6818
rect 20662 6778 20720 6784
rect 20854 6778 20912 6784
rect 21046 6778 21104 6784
rect 21238 6778 21296 6784
rect 21430 6778 21488 6784
rect 4091 6614 4149 6620
rect 4209 6614 4267 6620
rect 4327 6614 4385 6620
rect 4445 6614 4503 6620
rect 4563 6614 4621 6620
rect 4681 6614 4739 6620
rect 4799 6614 4857 6620
rect 4917 6614 4975 6620
rect 5035 6614 5093 6620
rect 5153 6614 5211 6620
rect 5599 6614 5657 6620
rect 5717 6614 5775 6620
rect 5835 6614 5893 6620
rect 5953 6614 6011 6620
rect 6071 6614 6129 6620
rect 6189 6614 6247 6620
rect 6307 6614 6365 6620
rect 6425 6614 6483 6620
rect 6543 6614 6601 6620
rect 6661 6614 6719 6620
rect 4091 6580 4103 6614
rect 4209 6580 4221 6614
rect 4327 6580 4339 6614
rect 4445 6580 4457 6614
rect 4563 6580 4575 6614
rect 4681 6580 4693 6614
rect 4799 6580 4811 6614
rect 4917 6580 4929 6614
rect 5035 6580 5047 6614
rect 5153 6580 5165 6614
rect 5599 6580 5611 6614
rect 5717 6580 5729 6614
rect 5835 6580 5847 6614
rect 5953 6580 5965 6614
rect 6071 6580 6083 6614
rect 6189 6580 6201 6614
rect 6307 6580 6319 6614
rect 6425 6580 6437 6614
rect 6543 6580 6555 6614
rect 6661 6580 6673 6614
rect 4091 6574 4149 6580
rect 4209 6574 4267 6580
rect 4327 6574 4385 6580
rect 4445 6574 4503 6580
rect 4563 6574 4621 6580
rect 4681 6574 4739 6580
rect 4799 6574 4857 6580
rect 4917 6574 4975 6580
rect 5035 6574 5093 6580
rect 5153 6574 5211 6580
rect 5599 6574 5657 6580
rect 5717 6574 5775 6580
rect 5835 6574 5893 6580
rect 5953 6574 6011 6580
rect 6071 6574 6129 6580
rect 6189 6574 6247 6580
rect 6307 6574 6365 6580
rect 6425 6574 6483 6580
rect 6543 6574 6601 6580
rect 6661 6574 6719 6580
rect 4091 6506 4149 6512
rect 4209 6506 4267 6512
rect 4327 6506 4385 6512
rect 4445 6506 4503 6512
rect 4563 6506 4621 6512
rect 4681 6506 4739 6512
rect 4799 6506 4857 6512
rect 4917 6506 4975 6512
rect 5035 6506 5093 6512
rect 5153 6506 5211 6512
rect 5599 6506 5657 6512
rect 5717 6506 5775 6512
rect 5835 6506 5893 6512
rect 5953 6506 6011 6512
rect 6071 6506 6129 6512
rect 6189 6506 6247 6512
rect 6307 6506 6365 6512
rect 6425 6506 6483 6512
rect 6543 6506 6601 6512
rect 6661 6506 6719 6512
rect 4091 6472 4103 6506
rect 4209 6472 4221 6506
rect 4327 6472 4339 6506
rect 4445 6472 4457 6506
rect 4563 6472 4575 6506
rect 4681 6472 4693 6506
rect 4799 6472 4811 6506
rect 4917 6472 4929 6506
rect 5035 6472 5047 6506
rect 5153 6472 5165 6506
rect 5599 6472 5611 6506
rect 5717 6472 5729 6506
rect 5835 6472 5847 6506
rect 5953 6472 5965 6506
rect 6071 6472 6083 6506
rect 6189 6472 6201 6506
rect 6307 6472 6319 6506
rect 6425 6472 6437 6506
rect 6543 6472 6555 6506
rect 6661 6472 6673 6506
rect 4091 6466 4149 6472
rect 4209 6466 4267 6472
rect 4327 6466 4385 6472
rect 4445 6466 4503 6472
rect 4563 6466 4621 6472
rect 4681 6466 4739 6472
rect 4799 6466 4857 6472
rect 4917 6466 4975 6472
rect 5035 6466 5093 6472
rect 5153 6466 5211 6472
rect 5599 6466 5657 6472
rect 5717 6466 5775 6472
rect 5835 6466 5893 6472
rect 5953 6466 6011 6472
rect 6071 6466 6129 6472
rect 6189 6466 6247 6472
rect 6307 6466 6365 6472
rect 6425 6466 6483 6472
rect 6543 6466 6601 6472
rect 6661 6466 6719 6472
rect 4091 6196 4149 6202
rect 4209 6196 4267 6202
rect 4327 6196 4385 6202
rect 4445 6196 4503 6202
rect 4563 6196 4621 6202
rect 4681 6196 4739 6202
rect 4799 6196 4857 6202
rect 4917 6196 4975 6202
rect 5035 6196 5093 6202
rect 5153 6196 5211 6202
rect 5599 6196 5657 6202
rect 5717 6196 5775 6202
rect 5835 6196 5893 6202
rect 5953 6196 6011 6202
rect 6071 6196 6129 6202
rect 6189 6196 6247 6202
rect 6307 6196 6365 6202
rect 6425 6196 6483 6202
rect 6543 6196 6601 6202
rect 6661 6196 6719 6202
rect 4091 6162 4103 6196
rect 4209 6162 4221 6196
rect 4327 6162 4339 6196
rect 4445 6162 4457 6196
rect 4563 6162 4575 6196
rect 4681 6162 4693 6196
rect 4799 6162 4811 6196
rect 4917 6162 4929 6196
rect 5035 6162 5047 6196
rect 5153 6162 5165 6196
rect 5599 6162 5611 6196
rect 5717 6162 5729 6196
rect 5835 6162 5847 6196
rect 5953 6162 5965 6196
rect 6071 6162 6083 6196
rect 6189 6162 6201 6196
rect 6307 6162 6319 6196
rect 6425 6162 6437 6196
rect 6543 6162 6555 6196
rect 6661 6162 6673 6196
rect 20650 6178 20708 6184
rect 20842 6178 20900 6184
rect 21034 6178 21092 6184
rect 21226 6178 21284 6184
rect 21418 6178 21476 6184
rect 4091 6156 4149 6162
rect 4209 6156 4267 6162
rect 4327 6156 4385 6162
rect 4445 6156 4503 6162
rect 4563 6156 4621 6162
rect 4681 6156 4739 6162
rect 4799 6156 4857 6162
rect 4917 6156 4975 6162
rect 5035 6156 5093 6162
rect 5153 6156 5211 6162
rect 5599 6156 5657 6162
rect 5717 6156 5775 6162
rect 5835 6156 5893 6162
rect 5953 6156 6011 6162
rect 6071 6156 6129 6162
rect 6189 6156 6247 6162
rect 6307 6156 6365 6162
rect 6425 6156 6483 6162
rect 6543 6156 6601 6162
rect 6661 6156 6719 6162
rect 20650 6144 20662 6178
rect 20842 6144 20854 6178
rect 21034 6144 21046 6178
rect 21226 6144 21238 6178
rect 21418 6144 21430 6178
rect 20650 6138 20708 6144
rect 20842 6138 20900 6144
rect 21034 6138 21092 6144
rect 21226 6138 21284 6144
rect 21418 6138 21476 6144
rect 4091 6088 4149 6094
rect 4209 6088 4267 6094
rect 4327 6088 4385 6094
rect 4445 6088 4503 6094
rect 4563 6088 4621 6094
rect 4681 6088 4739 6094
rect 4799 6088 4857 6094
rect 4917 6088 4975 6094
rect 5035 6088 5093 6094
rect 5153 6088 5211 6094
rect 5599 6088 5657 6094
rect 5717 6088 5775 6094
rect 5835 6088 5893 6094
rect 5953 6088 6011 6094
rect 6071 6088 6129 6094
rect 6189 6088 6247 6094
rect 6307 6088 6365 6094
rect 6425 6088 6483 6094
rect 6543 6088 6601 6094
rect 6661 6088 6719 6094
rect 4091 6054 4103 6088
rect 4209 6054 4221 6088
rect 4327 6054 4339 6088
rect 4445 6054 4457 6088
rect 4563 6054 4575 6088
rect 4681 6054 4693 6088
rect 4799 6054 4811 6088
rect 4917 6054 4929 6088
rect 5035 6054 5047 6088
rect 5153 6054 5165 6088
rect 5599 6054 5611 6088
rect 5717 6054 5729 6088
rect 5835 6054 5847 6088
rect 5953 6054 5965 6088
rect 6071 6054 6083 6088
rect 6189 6054 6201 6088
rect 6307 6054 6319 6088
rect 6425 6054 6437 6088
rect 6543 6054 6555 6088
rect 6661 6054 6673 6088
rect 4091 6048 4149 6054
rect 4209 6048 4267 6054
rect 4327 6048 4385 6054
rect 4445 6048 4503 6054
rect 4563 6048 4621 6054
rect 4681 6048 4739 6054
rect 4799 6048 4857 6054
rect 4917 6048 4975 6054
rect 5035 6048 5093 6054
rect 5153 6048 5211 6054
rect 5599 6048 5657 6054
rect 5717 6048 5775 6054
rect 5835 6048 5893 6054
rect 5953 6048 6011 6054
rect 6071 6048 6129 6054
rect 6189 6048 6247 6054
rect 6307 6048 6365 6054
rect 6425 6048 6483 6054
rect 6543 6048 6601 6054
rect 6661 6048 6719 6054
rect 4091 5778 4149 5784
rect 4209 5778 4267 5784
rect 4327 5778 4385 5784
rect 4445 5778 4503 5784
rect 4563 5778 4621 5784
rect 4681 5778 4739 5784
rect 4799 5778 4857 5784
rect 4917 5778 4975 5784
rect 5035 5778 5093 5784
rect 5153 5778 5211 5784
rect 5599 5778 5657 5784
rect 5717 5778 5775 5784
rect 5835 5778 5893 5784
rect 5953 5778 6011 5784
rect 6071 5778 6129 5784
rect 6189 5778 6247 5784
rect 6307 5778 6365 5784
rect 6425 5778 6483 5784
rect 6543 5778 6601 5784
rect 6661 5778 6719 5784
rect 4091 5744 4103 5778
rect 4209 5744 4221 5778
rect 4327 5744 4339 5778
rect 4445 5744 4457 5778
rect 4563 5744 4575 5778
rect 4681 5744 4693 5778
rect 4799 5744 4811 5778
rect 4917 5744 4929 5778
rect 5035 5744 5047 5778
rect 5153 5744 5165 5778
rect 5599 5744 5611 5778
rect 5717 5744 5729 5778
rect 5835 5744 5847 5778
rect 5953 5744 5965 5778
rect 6071 5744 6083 5778
rect 6189 5744 6201 5778
rect 6307 5744 6319 5778
rect 6425 5744 6437 5778
rect 6543 5744 6555 5778
rect 6661 5744 6673 5778
rect 4091 5738 4149 5744
rect 4209 5738 4267 5744
rect 4327 5738 4385 5744
rect 4445 5738 4503 5744
rect 4563 5738 4621 5744
rect 4681 5738 4739 5744
rect 4799 5738 4857 5744
rect 4917 5738 4975 5744
rect 5035 5738 5093 5744
rect 5153 5738 5211 5744
rect 5599 5738 5657 5744
rect 5717 5738 5775 5744
rect 5835 5738 5893 5744
rect 5953 5738 6011 5744
rect 6071 5738 6129 5744
rect 6189 5738 6247 5744
rect 6307 5738 6365 5744
rect 6425 5738 6483 5744
rect 6543 5738 6601 5744
rect 6661 5738 6719 5744
rect 20746 5268 20804 5274
rect 20938 5268 20996 5274
rect 21130 5268 21188 5274
rect 21322 5268 21380 5274
rect 21514 5268 21572 5274
rect 20746 5234 20758 5268
rect 20938 5234 20950 5268
rect 21130 5234 21142 5268
rect 21322 5234 21334 5268
rect 21514 5234 21526 5268
rect 20746 5228 20804 5234
rect 20938 5228 20996 5234
rect 21130 5228 21188 5234
rect 21322 5228 21380 5234
rect 21514 5228 21572 5234
rect 20746 5160 20804 5166
rect 20938 5160 20996 5166
rect 21130 5160 21188 5166
rect 21322 5160 21380 5166
rect 21514 5160 21572 5166
rect 20746 5126 20758 5160
rect 20938 5126 20950 5160
rect 21130 5126 21142 5160
rect 21322 5126 21334 5160
rect 21514 5126 21526 5160
rect 20746 5120 20804 5126
rect 20938 5120 20996 5126
rect 21130 5120 21188 5126
rect 21322 5120 21380 5126
rect 21514 5120 21572 5126
rect 20650 4250 20708 4256
rect 20842 4250 20900 4256
rect 21034 4250 21092 4256
rect 21226 4250 21284 4256
rect 21418 4250 21476 4256
rect 20650 4216 20662 4250
rect 20842 4216 20854 4250
rect 21034 4216 21046 4250
rect 21226 4216 21238 4250
rect 21418 4216 21430 4250
rect 20650 4210 20708 4216
rect 20842 4210 20900 4216
rect 21034 4210 21092 4216
rect 21226 4210 21284 4216
rect 21418 4210 21476 4216
rect 7987 3874 8045 3880
rect 8105 3874 8163 3880
rect 8223 3874 8281 3880
rect 8341 3874 8399 3880
rect 8459 3874 8517 3880
rect 8577 3874 8635 3880
rect 8695 3874 8753 3880
rect 8813 3874 8871 3880
rect 8931 3874 8989 3880
rect 9049 3874 9107 3880
rect 9167 3874 9225 3880
rect 9285 3874 9343 3880
rect 9403 3874 9461 3880
rect 9521 3874 9579 3880
rect 9639 3874 9697 3880
rect 9757 3874 9815 3880
rect 9875 3874 9933 3880
rect 9993 3874 10051 3880
rect 10111 3874 10169 3880
rect 10229 3874 10287 3880
rect 7987 3840 7999 3874
rect 8105 3840 8117 3874
rect 8223 3840 8235 3874
rect 8341 3840 8353 3874
rect 8459 3840 8471 3874
rect 8577 3840 8589 3874
rect 8695 3840 8707 3874
rect 8813 3840 8825 3874
rect 8931 3840 8943 3874
rect 9049 3840 9061 3874
rect 9167 3840 9179 3874
rect 9285 3840 9297 3874
rect 9403 3840 9415 3874
rect 9521 3840 9533 3874
rect 9639 3840 9651 3874
rect 9757 3840 9769 3874
rect 9875 3840 9887 3874
rect 9993 3840 10005 3874
rect 10111 3840 10123 3874
rect 10229 3840 10241 3874
rect 7987 3834 8045 3840
rect 8105 3834 8163 3840
rect 8223 3834 8281 3840
rect 8341 3834 8399 3840
rect 8459 3834 8517 3840
rect 8577 3834 8635 3840
rect 8695 3834 8753 3840
rect 8813 3834 8871 3840
rect 8931 3834 8989 3840
rect 9049 3834 9107 3840
rect 9167 3834 9225 3840
rect 9285 3834 9343 3840
rect 9403 3834 9461 3840
rect 9521 3834 9579 3840
rect 9639 3834 9697 3840
rect 9757 3834 9815 3840
rect 9875 3834 9933 3840
rect 9993 3834 10051 3840
rect 10111 3834 10169 3840
rect 10229 3834 10287 3840
rect 7987 3364 8045 3370
rect 8105 3364 8163 3370
rect 8223 3364 8281 3370
rect 8341 3364 8399 3370
rect 8459 3364 8517 3370
rect 8577 3364 8635 3370
rect 8695 3364 8753 3370
rect 8813 3364 8871 3370
rect 8931 3364 8989 3370
rect 9049 3364 9107 3370
rect 9167 3364 9225 3370
rect 9285 3364 9343 3370
rect 9403 3364 9461 3370
rect 9521 3364 9579 3370
rect 9639 3364 9697 3370
rect 9757 3364 9815 3370
rect 9875 3364 9933 3370
rect 9993 3364 10051 3370
rect 10111 3364 10169 3370
rect 10229 3364 10287 3370
rect 7987 3330 7999 3364
rect 8105 3330 8117 3364
rect 8223 3330 8235 3364
rect 8341 3330 8353 3364
rect 8459 3330 8471 3364
rect 8577 3330 8589 3364
rect 8695 3330 8707 3364
rect 8813 3330 8825 3364
rect 8931 3330 8943 3364
rect 9049 3330 9061 3364
rect 9167 3330 9179 3364
rect 9285 3330 9297 3364
rect 9403 3330 9415 3364
rect 9521 3330 9533 3364
rect 9639 3330 9651 3364
rect 9757 3330 9769 3364
rect 9875 3330 9887 3364
rect 9993 3330 10005 3364
rect 10111 3330 10123 3364
rect 10229 3330 10241 3364
rect 7987 3324 8045 3330
rect 8105 3324 8163 3330
rect 8223 3324 8281 3330
rect 8341 3324 8399 3330
rect 8459 3324 8517 3330
rect 8577 3324 8635 3330
rect 8695 3324 8753 3330
rect 8813 3324 8871 3330
rect 8931 3324 8989 3330
rect 9049 3324 9107 3330
rect 9167 3324 9225 3330
rect 9285 3324 9343 3330
rect 9403 3324 9461 3330
rect 9521 3324 9579 3330
rect 9639 3324 9697 3330
rect 9757 3324 9815 3330
rect 9875 3324 9933 3330
rect 9993 3324 10051 3330
rect 10111 3324 10169 3330
rect 10229 3324 10287 3330
<< pwell >>
rect 1872 7070 1982 7542
rect 2684 7472 2800 7944
<< viali >>
rect 4352 9918 4562 9988
rect 6330 9916 6522 9984
rect 8164 9936 8432 10006
rect 12314 9934 12618 10008
rect 14222 9936 14510 10006
rect 18376 9932 18668 10008
rect 20274 9878 20448 9954
rect 21366 9880 21528 9956
rect 1068 3292 1142 3556
rect 2038 2042 2246 2134
rect 4814 2046 5046 2134
rect 7516 2052 7754 2138
rect 10260 2052 10500 2136
rect 12758 2052 12986 2138
rect 15548 2054 15776 2136
rect 17912 2060 18164 2136
rect 20726 2056 20964 2136
<< metal1 >>
rect 30 10348 22606 10794
rect 102 8284 302 8484
rect 546 4831 752 10348
rect 4312 9988 4604 10348
rect 4312 9918 4352 9988
rect 4562 9918 4604 9988
rect 4312 9908 4604 9918
rect 6276 9984 6568 10348
rect 6276 9916 6330 9984
rect 6522 9916 6568 9984
rect 8088 10006 8492 10348
rect 8088 9936 8164 10006
rect 8432 9936 8492 10006
rect 8088 9922 8492 9936
rect 12264 10008 12668 10348
rect 12264 9934 12314 10008
rect 12618 9934 12668 10008
rect 12264 9920 12668 9934
rect 14158 10006 14562 10348
rect 14158 9936 14222 10006
rect 14510 9936 14562 10006
rect 14158 9924 14562 9936
rect 18324 10008 18728 10348
rect 18324 9932 18376 10008
rect 18668 9932 18728 10008
rect 18324 9922 18728 9932
rect 20240 9954 20478 10348
rect 6276 9906 6568 9916
rect 20240 9878 20274 9954
rect 20448 9878 20478 9954
rect 20240 9870 20478 9878
rect 21332 9956 21570 10348
rect 21332 9880 21366 9956
rect 21528 9880 21570 9956
rect 21332 9866 21570 9880
rect 2293 7542 2403 7941
rect 1128 7436 1610 7536
rect 1128 7074 1222 7436
rect 1510 7080 1610 7436
rect 1872 7432 2403 7542
rect 2684 7828 3202 7944
rect 2684 7472 2800 7828
rect 3086 7450 3202 7828
rect 1872 7070 1982 7432
rect 22378 6402 22578 6602
rect 1113 4831 1238 5454
rect 1502 5172 1606 5528
rect 1878 5172 1982 5524
rect 1502 5068 1982 5172
rect 2290 5178 2404 5528
rect 2689 5178 2803 5549
rect 2290 5064 2803 5178
rect 546 4632 1240 4831
rect 22380 4698 22580 4898
rect 98 4186 298 4386
rect 1218 3627 6304 3630
rect 516 3556 1148 3582
rect 1218 3556 6569 3627
rect 516 3292 1068 3556
rect 1142 3292 1148 3556
rect 6255 3553 6569 3556
rect 1190 3460 1200 3522
rect 1256 3460 1266 3522
rect 2106 3460 2116 3522
rect 2172 3460 2182 3522
rect 3022 3460 3032 3522
rect 3088 3460 3098 3522
rect 3938 3460 3948 3522
rect 4004 3460 4014 3522
rect 4852 3456 4862 3518
rect 4918 3456 4928 3518
rect 5768 3458 5778 3520
rect 5834 3458 5844 3520
rect 1642 3318 1652 3374
rect 1722 3318 1732 3374
rect 2558 3318 2568 3374
rect 2638 3318 2648 3374
rect 3472 3320 3482 3376
rect 3552 3320 3562 3376
rect 4390 3318 4400 3374
rect 4470 3318 4480 3374
rect 5306 3318 5316 3374
rect 5386 3318 5396 3374
rect 516 3272 1148 3292
rect 6495 3282 6569 3553
rect 575 1536 768 3272
rect 1222 3208 6569 3282
rect 1972 2134 2310 2148
rect 1972 2042 2038 2134
rect 2246 2042 2310 2134
rect 575 1528 830 1536
rect 1972 1528 2310 2042
rect 4762 2134 5098 2148
rect 4762 2046 4814 2134
rect 5046 2046 5098 2134
rect 4762 1528 5098 2046
rect 7462 2138 7800 2150
rect 7462 2052 7516 2138
rect 7754 2052 7800 2138
rect 7462 1528 7800 2052
rect 10206 2136 10546 2148
rect 10206 2052 10260 2136
rect 10500 2052 10546 2136
rect 10206 1528 10546 2052
rect 12692 2138 13036 2150
rect 12692 2052 12758 2138
rect 12986 2052 13036 2138
rect 12692 1528 13036 2052
rect 15488 2136 15834 2148
rect 15488 2054 15548 2136
rect 15776 2054 15834 2136
rect 15488 1528 15834 2054
rect 17864 2136 18210 2148
rect 17864 2060 17912 2136
rect 18164 2060 18210 2136
rect 17864 2052 18210 2060
rect 20676 2136 21024 2148
rect 20676 2056 20726 2136
rect 20964 2056 21024 2136
rect 17864 1528 18212 2052
rect 20676 1528 21024 2056
rect 10 1082 22586 1528
rect 17864 1078 18212 1082
<< via1 >>
rect 1200 3460 1256 3522
rect 2116 3460 2172 3522
rect 3032 3460 3088 3522
rect 3948 3460 4004 3522
rect 4862 3456 4918 3518
rect 5778 3458 5834 3520
rect 1652 3318 1722 3374
rect 2568 3318 2638 3374
rect 3482 3320 3552 3376
rect 4400 3318 4470 3374
rect 5316 3318 5386 3374
<< metal2 >>
rect 1200 3522 1256 3532
rect 2116 3522 2172 3532
rect 3032 3522 3088 3532
rect 3948 3522 4004 3532
rect 4862 3522 4918 3528
rect 5778 3522 5834 3530
rect 1182 3460 1200 3522
rect 1256 3460 2116 3522
rect 2172 3460 3032 3522
rect 3088 3460 3948 3522
rect 4004 3520 6200 3522
rect 4004 3518 5778 3520
rect 4004 3460 4862 3518
rect 1182 3458 4862 3460
rect 1200 3450 1256 3458
rect 2116 3450 2172 3458
rect 3032 3450 3088 3458
rect 3948 3450 4004 3458
rect 4918 3458 5778 3518
rect 5834 3458 6200 3520
rect 4862 3446 4918 3456
rect 5778 3448 5834 3458
rect 1652 3374 1722 3384
rect 2568 3374 2638 3384
rect 3482 3376 3552 3386
rect 1180 3318 1652 3374
rect 1722 3318 2568 3374
rect 2638 3320 3482 3374
rect 4400 3374 4470 3384
rect 5316 3374 5386 3384
rect 3552 3320 4400 3374
rect 2638 3318 4400 3320
rect 4470 3318 5316 3374
rect 5386 3318 6200 3374
rect 1180 3312 6200 3318
rect 1652 3308 1722 3312
rect 2568 3308 2638 3312
rect 3482 3310 3552 3312
rect 4400 3308 4470 3312
rect 5316 3308 5386 3312
use sky130_fd_pr__nfet_01v8_FMJ72H  XM1
timestamp 1713266475
transform 1 0 4651 0 1 6752
box -757 -1146 757 1146
use sky130_fd_pr__nfet_01v8_FMJ72H  XM2
timestamp 1713266475
transform 1 0 6159 0 1 6752
box -757 -1146 757 1146
use sky130_fd_pr__pfet_01v8_3H5TVM  XM3
timestamp 1713266475
transform 1 0 6410 0 1 9677
box -812 -319 812 319
use sky130_fd_pr__pfet_01v8_3H5TVM  XM4
timestamp 1713266475
transform 1 0 4454 0 1 9683
box -812 -319 812 319
use sky130_fd_pr__nfet_01v8_EPHDNF  XM5
timestamp 1713266475
transform 1 0 3517 0 1 3420
box -2457 -310 2457 310
use sky130_fd_pr__nfet_01v8_EPHDNF  XM6
timestamp 1713266475
transform 1 0 3517 0 1 2358
box -2457 -310 2457 310
use sky130_fd_pr__nfet_01v8_SMX62R  XM7
timestamp 1713266475
transform 1 0 9137 0 1 3602
box -1347 -410 1347 410
use sky130_fd_pr__nfet_01v8_EPHDNF  XM8
timestamp 1713266475
transform 1 0 8991 0 1 2356
box -2457 -310 2457 310
use sky130_fd_pr__pfet_01v8_P7N2DR  XM9
timestamp 1713266475
transform 1 0 10459 0 1 7343
box -2747 -2677 2747 2677
use sky130_fd_pr__pfet_01v8_P7N2DR  XM10
timestamp 1713266475
transform 1 0 16531 0 1 7343
box -2747 -2677 2747 2677
use sky130_fd_pr__nfet_01v8_EPHDNF  XM11
timestamp 1713266475
transform 1 0 14255 0 1 2358
box -2457 -310 2457 310
use sky130_fd_pr__nfet_01v8_V5FT3Q  XM12
timestamp 1713266475
transform 1 0 20546 0 1 3358
box -1312 -410 1312 410
use sky130_fd_pr__pfet_01v8_3HZ9VM  XM13
timestamp 1713266475
transform 1 0 20354 0 1 9245
box -296 -719 296 719
use sky130_fd_pr__nfet_01v8_EPHDNF  XM14
timestamp 1713266475
transform 1 0 19417 0 1 2358
box -2457 -310 2457 310
use sky130_fd_pr__nfet_01v8_GSBCLJ  XM15
timestamp 1713266475
transform 1 0 21111 0 1 5197
box -647 -1119 647 1119
use sky130_fd_pr__pfet_01v8_3HZ9VM  XM16
timestamp 1713266475
transform 1 0 21446 0 1 9243
box -296 -719 296 719
use sky130_fd_pr__pfet_01v8_BDVWJN  XM17
timestamp 1713266475
transform 1 0 21123 0 1 7365
box -647 -719 647 719
use sky130_fd_pr__res_xhigh_po_0p35_RF5GSL  XR1
timestamp 1713266475
transform 1 0 1553 0 1 6304
box -201 -1382 201 1382
use sky130_fd_pr__res_xhigh_po_0p35_RF5GSL  XR2
timestamp 1713266475
transform 1 0 1161 0 1 6304
box -201 -1382 201 1382
use sky130_fd_pr__res_xhigh_po_0p35_RF5GSL  XR3
timestamp 1713266475
transform 1 0 1945 0 1 6304
box -201 -1382 201 1382
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR4
timestamp 1713266475
transform 1 0 2345 0 1 6500
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR5
timestamp 1713266475
transform 1 0 3143 0 1 6500
box -201 -1582 201 1582
use sky130_fd_pr__res_high_po_0p35_FFK5MY  XR6
timestamp 1713266475
transform 1 0 2747 0 1 6510
box -201 -1582 201 1582
<< labels >>
flabel metal1 106 1246 306 1446 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 22378 6402 22578 6602 0 FreeSans 256 0 0 0 z
port 2 nsew
flabel metal1 22380 4698 22580 4898 0 FreeSans 256 0 0 0 x
port 5 nsew
flabel metal1 98 4186 298 4386 0 FreeSans 256 0 0 0 y
port 3 nsew
flabel metal1 102 8284 302 8484 0 FreeSans 256 0 0 0 ref
port 4 nsew
flabel metal1 92 10506 292 10706 0 FreeSans 256 0 0 0 vdd
port 0 nsew
<< end >>
