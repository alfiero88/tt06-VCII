** sch_path: /home/ttuser/tt06-VCII/xschem/VCII-testbench.sch
**.subckt VCII-testbench
V1 vdd GND 1.8
V2 GND vss 0
V3 Ref vss 0.9
x1 vdd vss net2 y Ref x VCII-final
I2 y Ref 0 ac 1 0 sin(0 2u 100K 0 0 0)
R1 x net1 10k m=1
Vmeas2 net1 Ref 0
.save i(vmeas2)
C1 net2 vss 5p m=1
R2 z net2 500 m=1
**** begin user architecture code



*save
*+ @m.xm1.msky130_fd_pr__nfet_01v8[gm]
*+ @m.xm2.msky130_fd_pr__nfet_01v8[gm]
*+ @m.xm4.msky130_fd_pr__pfet_01v8[gm]
*+ @m.xm3.msky130_fd_pr__pfet_01v8[gm]

.options savecurrents
.control
  save all
  op
  remzerovec
  write VCII-testbench.raw
  set appendwrite
  dc temp -40 140 1
  write VCII-testbench.raw
  ac dec 100 1 1e12
  remzerovec
  write VCII-testbench.raw
  tran 0.1n 10u
  write VCII-testbench.raw
  *quit 0
.endc




.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  VCII-final.sym # of pins=6
** sym_path: /home/ttuser/tt06-VCII/xschem/VCII-final.sym
** sch_path: /home/ttuser/tt06-VCII/xschem/VCII-final.sch
.subckt VCII-final vdd vss z y ref x
*.iopin x
*.iopin y
*.iopin z
*.iopin vdd
*.iopin vss
*.iopin ref
XM1 G1 ref B1 vss sky130_fd_pr__nfet_01v8 L=0.3 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM2 D1 y B1 vss sky130_fd_pr__nfet_01v8 L=0.3 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM3 D1 G1 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=5 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 G1 G1 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=5 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 B1 G2 vss vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 G2 G2 vss vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 G3 D1 y vss sky130_fd_pr__nfet_01v8 L=0.3 W=40 nf=20 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 y G2 vss vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 G3 G3 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=50 nf=20 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=7 m=7
XM10 x G3 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=50 nf=20 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=7 m=7
XM11 x G2 vss vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 net1 G2 vss vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 z G2 vss vss sky130_fd_pr__nfet_01v8 L=2 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 vdd G4 z vss sky130_fd_pr__nfet_01v8 L=0.15 W=40 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM13 net1 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 G4 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 vss x G4 vdd sky130_fd_pr__pfet_01v8 L=0.15 W=50 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR2 net2 vdd vss sky130_fd_pr__res_xhigh_po_0p35 L=8 mult=1 m=1
XR1 net3 net2 vss sky130_fd_pr__res_xhigh_po_0p35 L=8 mult=1 m=1
XR3 net4 net3 vss sky130_fd_pr__res_xhigh_po_0p35 L=8 mult=1 m=1
XR5 net6 net5 vss sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR6 net5 G2 vss sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR4 net4 net6 vss sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
.ends

.GLOBAL GND
.end
