** sch_path: /home/ttuser/tt06-VCII/xschem/VCII-final.sch
.subckt VCII-final vdd vss z y ref x
*.PININFO x:B y:B z:B vdd:B vss:B ref:B
XM1 G1 ref B1 vss sky130_fd_pr__nfet_01v8 L=0.3 W=10 nf=10 m=5
XM2 D1 y B1 vss sky130_fd_pr__nfet_01v8 L=0.3 W=10 nf=10 m=5
XM3 D1 G1 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=5 nf=5 m=1
XM4 G1 G1 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=5 nf=5 m=1
XM5 B1 G2 vss vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=10 m=1
XM6 G2 G2 vss vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=10 m=1
XM7 G3 D1 y vss sky130_fd_pr__nfet_01v8 L=0.3 W=40 nf=20 m=1
XM8 y G2 vss vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=10 m=1
XM9 G3 G3 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=50 nf=20 m=7
XM10 x G3 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=50 nf=20 m=7
XM11 x G2 vss vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=10 m=1
XM14 net1 G2 vss vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=10 m=1
XM12 z G2 vss vss sky130_fd_pr__nfet_01v8 L=2 W=2 nf=2 m=1
XM15 vdd G4 z vss sky130_fd_pr__nfet_01v8 L=0.15 W=40 nf=10 m=2
XM13 net1 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=5 nf=1 m=1
XM16 G4 net1 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=5 nf=1 m=1
XM17 vss x G4 vdd sky130_fd_pr__pfet_01v8 L=0.15 W=50 nf=10 m=1
XR2 net2 vdd vss sky130_fd_pr__res_xhigh_po_0p35 L=8 mult=1 m=1
XR1 net3 net2 vss sky130_fd_pr__res_xhigh_po_0p35 L=8 mult=1 m=1
XR3 net4 net3 vss sky130_fd_pr__res_xhigh_po_0p35 L=8 mult=1 m=1
XR5 net6 net5 vss sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR6 net5 G2 vss sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XR4 net4 net6 vss sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
.ends
.end
