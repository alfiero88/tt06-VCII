magic
tech sky130A
magscale 1 2
timestamp 1713266475
<< error_p >>
rect -560 1008 -502 1014
rect -442 1008 -384 1014
rect -324 1008 -266 1014
rect -206 1008 -148 1014
rect -88 1008 -30 1014
rect 30 1008 88 1014
rect 148 1008 206 1014
rect 266 1008 324 1014
rect 384 1008 442 1014
rect 502 1008 560 1014
rect -560 974 -548 1008
rect -442 974 -430 1008
rect -324 974 -312 1008
rect -206 974 -194 1008
rect -88 974 -76 1008
rect 30 974 42 1008
rect 148 974 160 1008
rect 266 974 278 1008
rect 384 974 396 1008
rect 502 974 514 1008
rect -560 968 -502 974
rect -442 968 -384 974
rect -324 968 -266 974
rect -206 968 -148 974
rect -88 968 -30 974
rect 30 968 88 974
rect 148 968 206 974
rect 266 968 324 974
rect 384 968 442 974
rect 502 968 560 974
rect -560 698 -502 704
rect -442 698 -384 704
rect -324 698 -266 704
rect -206 698 -148 704
rect -88 698 -30 704
rect 30 698 88 704
rect 148 698 206 704
rect 266 698 324 704
rect 384 698 442 704
rect 502 698 560 704
rect -560 664 -548 698
rect -442 664 -430 698
rect -324 664 -312 698
rect -206 664 -194 698
rect -88 664 -76 698
rect 30 664 42 698
rect 148 664 160 698
rect 266 664 278 698
rect 384 664 396 698
rect 502 664 514 698
rect -560 658 -502 664
rect -442 658 -384 664
rect -324 658 -266 664
rect -206 658 -148 664
rect -88 658 -30 664
rect 30 658 88 664
rect 148 658 206 664
rect 266 658 324 664
rect 384 658 442 664
rect 502 658 560 664
rect -560 590 -502 596
rect -442 590 -384 596
rect -324 590 -266 596
rect -206 590 -148 596
rect -88 590 -30 596
rect 30 590 88 596
rect 148 590 206 596
rect 266 590 324 596
rect 384 590 442 596
rect 502 590 560 596
rect -560 556 -548 590
rect -442 556 -430 590
rect -324 556 -312 590
rect -206 556 -194 590
rect -88 556 -76 590
rect 30 556 42 590
rect 148 556 160 590
rect 266 556 278 590
rect 384 556 396 590
rect 502 556 514 590
rect -560 550 -502 556
rect -442 550 -384 556
rect -324 550 -266 556
rect -206 550 -148 556
rect -88 550 -30 556
rect 30 550 88 556
rect 148 550 206 556
rect 266 550 324 556
rect 384 550 442 556
rect 502 550 560 556
rect -560 280 -502 286
rect -442 280 -384 286
rect -324 280 -266 286
rect -206 280 -148 286
rect -88 280 -30 286
rect 30 280 88 286
rect 148 280 206 286
rect 266 280 324 286
rect 384 280 442 286
rect 502 280 560 286
rect -560 246 -548 280
rect -442 246 -430 280
rect -324 246 -312 280
rect -206 246 -194 280
rect -88 246 -76 280
rect 30 246 42 280
rect 148 246 160 280
rect 266 246 278 280
rect 384 246 396 280
rect 502 246 514 280
rect -560 240 -502 246
rect -442 240 -384 246
rect -324 240 -266 246
rect -206 240 -148 246
rect -88 240 -30 246
rect 30 240 88 246
rect 148 240 206 246
rect 266 240 324 246
rect 384 240 442 246
rect 502 240 560 246
rect -560 172 -502 178
rect -442 172 -384 178
rect -324 172 -266 178
rect -206 172 -148 178
rect -88 172 -30 178
rect 30 172 88 178
rect 148 172 206 178
rect 266 172 324 178
rect 384 172 442 178
rect 502 172 560 178
rect -560 138 -548 172
rect -442 138 -430 172
rect -324 138 -312 172
rect -206 138 -194 172
rect -88 138 -76 172
rect 30 138 42 172
rect 148 138 160 172
rect 266 138 278 172
rect 384 138 396 172
rect 502 138 514 172
rect -560 132 -502 138
rect -442 132 -384 138
rect -324 132 -266 138
rect -206 132 -148 138
rect -88 132 -30 138
rect 30 132 88 138
rect 148 132 206 138
rect 266 132 324 138
rect 384 132 442 138
rect 502 132 560 138
rect -560 -138 -502 -132
rect -442 -138 -384 -132
rect -324 -138 -266 -132
rect -206 -138 -148 -132
rect -88 -138 -30 -132
rect 30 -138 88 -132
rect 148 -138 206 -132
rect 266 -138 324 -132
rect 384 -138 442 -132
rect 502 -138 560 -132
rect -560 -172 -548 -138
rect -442 -172 -430 -138
rect -324 -172 -312 -138
rect -206 -172 -194 -138
rect -88 -172 -76 -138
rect 30 -172 42 -138
rect 148 -172 160 -138
rect 266 -172 278 -138
rect 384 -172 396 -138
rect 502 -172 514 -138
rect -560 -178 -502 -172
rect -442 -178 -384 -172
rect -324 -178 -266 -172
rect -206 -178 -148 -172
rect -88 -178 -30 -172
rect 30 -178 88 -172
rect 148 -178 206 -172
rect 266 -178 324 -172
rect 384 -178 442 -172
rect 502 -178 560 -172
rect -560 -246 -502 -240
rect -442 -246 -384 -240
rect -324 -246 -266 -240
rect -206 -246 -148 -240
rect -88 -246 -30 -240
rect 30 -246 88 -240
rect 148 -246 206 -240
rect 266 -246 324 -240
rect 384 -246 442 -240
rect 502 -246 560 -240
rect -560 -280 -548 -246
rect -442 -280 -430 -246
rect -324 -280 -312 -246
rect -206 -280 -194 -246
rect -88 -280 -76 -246
rect 30 -280 42 -246
rect 148 -280 160 -246
rect 266 -280 278 -246
rect 384 -280 396 -246
rect 502 -280 514 -246
rect -560 -286 -502 -280
rect -442 -286 -384 -280
rect -324 -286 -266 -280
rect -206 -286 -148 -280
rect -88 -286 -30 -280
rect 30 -286 88 -280
rect 148 -286 206 -280
rect 266 -286 324 -280
rect 384 -286 442 -280
rect 502 -286 560 -280
rect -560 -556 -502 -550
rect -442 -556 -384 -550
rect -324 -556 -266 -550
rect -206 -556 -148 -550
rect -88 -556 -30 -550
rect 30 -556 88 -550
rect 148 -556 206 -550
rect 266 -556 324 -550
rect 384 -556 442 -550
rect 502 -556 560 -550
rect -560 -590 -548 -556
rect -442 -590 -430 -556
rect -324 -590 -312 -556
rect -206 -590 -194 -556
rect -88 -590 -76 -556
rect 30 -590 42 -556
rect 148 -590 160 -556
rect 266 -590 278 -556
rect 384 -590 396 -556
rect 502 -590 514 -556
rect -560 -596 -502 -590
rect -442 -596 -384 -590
rect -324 -596 -266 -590
rect -206 -596 -148 -590
rect -88 -596 -30 -590
rect 30 -596 88 -590
rect 148 -596 206 -590
rect 266 -596 324 -590
rect 384 -596 442 -590
rect 502 -596 560 -590
rect -560 -664 -502 -658
rect -442 -664 -384 -658
rect -324 -664 -266 -658
rect -206 -664 -148 -658
rect -88 -664 -30 -658
rect 30 -664 88 -658
rect 148 -664 206 -658
rect 266 -664 324 -658
rect 384 -664 442 -658
rect 502 -664 560 -658
rect -560 -698 -548 -664
rect -442 -698 -430 -664
rect -324 -698 -312 -664
rect -206 -698 -194 -664
rect -88 -698 -76 -664
rect 30 -698 42 -664
rect 148 -698 160 -664
rect 266 -698 278 -664
rect 384 -698 396 -664
rect 502 -698 514 -664
rect -560 -704 -502 -698
rect -442 -704 -384 -698
rect -324 -704 -266 -698
rect -206 -704 -148 -698
rect -88 -704 -30 -698
rect 30 -704 88 -698
rect 148 -704 206 -698
rect 266 -704 324 -698
rect 384 -704 442 -698
rect 502 -704 560 -698
rect -560 -974 -502 -968
rect -442 -974 -384 -968
rect -324 -974 -266 -968
rect -206 -974 -148 -968
rect -88 -974 -30 -968
rect 30 -974 88 -968
rect 148 -974 206 -968
rect 266 -974 324 -968
rect 384 -974 442 -968
rect 502 -974 560 -968
rect -560 -1008 -548 -974
rect -442 -1008 -430 -974
rect -324 -1008 -312 -974
rect -206 -1008 -194 -974
rect -88 -1008 -76 -974
rect 30 -1008 42 -974
rect 148 -1008 160 -974
rect 266 -1008 278 -974
rect 384 -1008 396 -974
rect 502 -1008 514 -974
rect -560 -1014 -502 -1008
rect -442 -1014 -384 -1008
rect -324 -1014 -266 -1008
rect -206 -1014 -148 -1008
rect -88 -1014 -30 -1008
rect 30 -1014 88 -1008
rect 148 -1014 206 -1008
rect 266 -1014 324 -1008
rect 384 -1014 442 -1008
rect 502 -1014 560 -1008
<< pwell >>
rect -757 -1146 757 1146
<< nmos >>
rect -561 736 -501 936
rect -443 736 -383 936
rect -325 736 -265 936
rect -207 736 -147 936
rect -89 736 -29 936
rect 29 736 89 936
rect 147 736 207 936
rect 265 736 325 936
rect 383 736 443 936
rect 501 736 561 936
rect -561 318 -501 518
rect -443 318 -383 518
rect -325 318 -265 518
rect -207 318 -147 518
rect -89 318 -29 518
rect 29 318 89 518
rect 147 318 207 518
rect 265 318 325 518
rect 383 318 443 518
rect 501 318 561 518
rect -561 -100 -501 100
rect -443 -100 -383 100
rect -325 -100 -265 100
rect -207 -100 -147 100
rect -89 -100 -29 100
rect 29 -100 89 100
rect 147 -100 207 100
rect 265 -100 325 100
rect 383 -100 443 100
rect 501 -100 561 100
rect -561 -518 -501 -318
rect -443 -518 -383 -318
rect -325 -518 -265 -318
rect -207 -518 -147 -318
rect -89 -518 -29 -318
rect 29 -518 89 -318
rect 147 -518 207 -318
rect 265 -518 325 -318
rect 383 -518 443 -318
rect 501 -518 561 -318
rect -561 -936 -501 -736
rect -443 -936 -383 -736
rect -325 -936 -265 -736
rect -207 -936 -147 -736
rect -89 -936 -29 -736
rect 29 -936 89 -736
rect 147 -936 207 -736
rect 265 -936 325 -736
rect 383 -936 443 -736
rect 501 -936 561 -736
<< ndiff >>
rect -619 924 -561 936
rect -619 748 -607 924
rect -573 748 -561 924
rect -619 736 -561 748
rect -501 924 -443 936
rect -501 748 -489 924
rect -455 748 -443 924
rect -501 736 -443 748
rect -383 924 -325 936
rect -383 748 -371 924
rect -337 748 -325 924
rect -383 736 -325 748
rect -265 924 -207 936
rect -265 748 -253 924
rect -219 748 -207 924
rect -265 736 -207 748
rect -147 924 -89 936
rect -147 748 -135 924
rect -101 748 -89 924
rect -147 736 -89 748
rect -29 924 29 936
rect -29 748 -17 924
rect 17 748 29 924
rect -29 736 29 748
rect 89 924 147 936
rect 89 748 101 924
rect 135 748 147 924
rect 89 736 147 748
rect 207 924 265 936
rect 207 748 219 924
rect 253 748 265 924
rect 207 736 265 748
rect 325 924 383 936
rect 325 748 337 924
rect 371 748 383 924
rect 325 736 383 748
rect 443 924 501 936
rect 443 748 455 924
rect 489 748 501 924
rect 443 736 501 748
rect 561 924 619 936
rect 561 748 573 924
rect 607 748 619 924
rect 561 736 619 748
rect -619 506 -561 518
rect -619 330 -607 506
rect -573 330 -561 506
rect -619 318 -561 330
rect -501 506 -443 518
rect -501 330 -489 506
rect -455 330 -443 506
rect -501 318 -443 330
rect -383 506 -325 518
rect -383 330 -371 506
rect -337 330 -325 506
rect -383 318 -325 330
rect -265 506 -207 518
rect -265 330 -253 506
rect -219 330 -207 506
rect -265 318 -207 330
rect -147 506 -89 518
rect -147 330 -135 506
rect -101 330 -89 506
rect -147 318 -89 330
rect -29 506 29 518
rect -29 330 -17 506
rect 17 330 29 506
rect -29 318 29 330
rect 89 506 147 518
rect 89 330 101 506
rect 135 330 147 506
rect 89 318 147 330
rect 207 506 265 518
rect 207 330 219 506
rect 253 330 265 506
rect 207 318 265 330
rect 325 506 383 518
rect 325 330 337 506
rect 371 330 383 506
rect 325 318 383 330
rect 443 506 501 518
rect 443 330 455 506
rect 489 330 501 506
rect 443 318 501 330
rect 561 506 619 518
rect 561 330 573 506
rect 607 330 619 506
rect 561 318 619 330
rect -619 88 -561 100
rect -619 -88 -607 88
rect -573 -88 -561 88
rect -619 -100 -561 -88
rect -501 88 -443 100
rect -501 -88 -489 88
rect -455 -88 -443 88
rect -501 -100 -443 -88
rect -383 88 -325 100
rect -383 -88 -371 88
rect -337 -88 -325 88
rect -383 -100 -325 -88
rect -265 88 -207 100
rect -265 -88 -253 88
rect -219 -88 -207 88
rect -265 -100 -207 -88
rect -147 88 -89 100
rect -147 -88 -135 88
rect -101 -88 -89 88
rect -147 -100 -89 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 89 88 147 100
rect 89 -88 101 88
rect 135 -88 147 88
rect 89 -100 147 -88
rect 207 88 265 100
rect 207 -88 219 88
rect 253 -88 265 88
rect 207 -100 265 -88
rect 325 88 383 100
rect 325 -88 337 88
rect 371 -88 383 88
rect 325 -100 383 -88
rect 443 88 501 100
rect 443 -88 455 88
rect 489 -88 501 88
rect 443 -100 501 -88
rect 561 88 619 100
rect 561 -88 573 88
rect 607 -88 619 88
rect 561 -100 619 -88
rect -619 -330 -561 -318
rect -619 -506 -607 -330
rect -573 -506 -561 -330
rect -619 -518 -561 -506
rect -501 -330 -443 -318
rect -501 -506 -489 -330
rect -455 -506 -443 -330
rect -501 -518 -443 -506
rect -383 -330 -325 -318
rect -383 -506 -371 -330
rect -337 -506 -325 -330
rect -383 -518 -325 -506
rect -265 -330 -207 -318
rect -265 -506 -253 -330
rect -219 -506 -207 -330
rect -265 -518 -207 -506
rect -147 -330 -89 -318
rect -147 -506 -135 -330
rect -101 -506 -89 -330
rect -147 -518 -89 -506
rect -29 -330 29 -318
rect -29 -506 -17 -330
rect 17 -506 29 -330
rect -29 -518 29 -506
rect 89 -330 147 -318
rect 89 -506 101 -330
rect 135 -506 147 -330
rect 89 -518 147 -506
rect 207 -330 265 -318
rect 207 -506 219 -330
rect 253 -506 265 -330
rect 207 -518 265 -506
rect 325 -330 383 -318
rect 325 -506 337 -330
rect 371 -506 383 -330
rect 325 -518 383 -506
rect 443 -330 501 -318
rect 443 -506 455 -330
rect 489 -506 501 -330
rect 443 -518 501 -506
rect 561 -330 619 -318
rect 561 -506 573 -330
rect 607 -506 619 -330
rect 561 -518 619 -506
rect -619 -748 -561 -736
rect -619 -924 -607 -748
rect -573 -924 -561 -748
rect -619 -936 -561 -924
rect -501 -748 -443 -736
rect -501 -924 -489 -748
rect -455 -924 -443 -748
rect -501 -936 -443 -924
rect -383 -748 -325 -736
rect -383 -924 -371 -748
rect -337 -924 -325 -748
rect -383 -936 -325 -924
rect -265 -748 -207 -736
rect -265 -924 -253 -748
rect -219 -924 -207 -748
rect -265 -936 -207 -924
rect -147 -748 -89 -736
rect -147 -924 -135 -748
rect -101 -924 -89 -748
rect -147 -936 -89 -924
rect -29 -748 29 -736
rect -29 -924 -17 -748
rect 17 -924 29 -748
rect -29 -936 29 -924
rect 89 -748 147 -736
rect 89 -924 101 -748
rect 135 -924 147 -748
rect 89 -936 147 -924
rect 207 -748 265 -736
rect 207 -924 219 -748
rect 253 -924 265 -748
rect 207 -936 265 -924
rect 325 -748 383 -736
rect 325 -924 337 -748
rect 371 -924 383 -748
rect 325 -936 383 -924
rect 443 -748 501 -736
rect 443 -924 455 -748
rect 489 -924 501 -748
rect 443 -936 501 -924
rect 561 -748 619 -736
rect 561 -924 573 -748
rect 607 -924 619 -748
rect 561 -936 619 -924
<< ndiffc >>
rect -607 748 -573 924
rect -489 748 -455 924
rect -371 748 -337 924
rect -253 748 -219 924
rect -135 748 -101 924
rect -17 748 17 924
rect 101 748 135 924
rect 219 748 253 924
rect 337 748 371 924
rect 455 748 489 924
rect 573 748 607 924
rect -607 330 -573 506
rect -489 330 -455 506
rect -371 330 -337 506
rect -253 330 -219 506
rect -135 330 -101 506
rect -17 330 17 506
rect 101 330 135 506
rect 219 330 253 506
rect 337 330 371 506
rect 455 330 489 506
rect 573 330 607 506
rect -607 -88 -573 88
rect -489 -88 -455 88
rect -371 -88 -337 88
rect -253 -88 -219 88
rect -135 -88 -101 88
rect -17 -88 17 88
rect 101 -88 135 88
rect 219 -88 253 88
rect 337 -88 371 88
rect 455 -88 489 88
rect 573 -88 607 88
rect -607 -506 -573 -330
rect -489 -506 -455 -330
rect -371 -506 -337 -330
rect -253 -506 -219 -330
rect -135 -506 -101 -330
rect -17 -506 17 -330
rect 101 -506 135 -330
rect 219 -506 253 -330
rect 337 -506 371 -330
rect 455 -506 489 -330
rect 573 -506 607 -330
rect -607 -924 -573 -748
rect -489 -924 -455 -748
rect -371 -924 -337 -748
rect -253 -924 -219 -748
rect -135 -924 -101 -748
rect -17 -924 17 -748
rect 101 -924 135 -748
rect 219 -924 253 -748
rect 337 -924 371 -748
rect 455 -924 489 -748
rect 573 -924 607 -748
<< psubdiff >>
rect -721 1076 -625 1110
rect 625 1076 721 1110
rect -721 1014 -687 1076
rect 687 1014 721 1076
rect -721 -1076 -687 -1014
rect 687 -1076 721 -1014
rect -721 -1110 -625 -1076
rect 625 -1110 721 -1076
<< psubdiffcont >>
rect -625 1076 625 1110
rect -721 -1014 -687 1014
rect 687 -1014 721 1014
rect -625 -1110 625 -1076
<< poly >>
rect -564 1008 -498 1024
rect -564 974 -548 1008
rect -514 974 -498 1008
rect -564 958 -498 974
rect -446 1008 -380 1024
rect -446 974 -430 1008
rect -396 974 -380 1008
rect -446 958 -380 974
rect -328 1008 -262 1024
rect -328 974 -312 1008
rect -278 974 -262 1008
rect -328 958 -262 974
rect -210 1008 -144 1024
rect -210 974 -194 1008
rect -160 974 -144 1008
rect -210 958 -144 974
rect -92 1008 -26 1024
rect -92 974 -76 1008
rect -42 974 -26 1008
rect -92 958 -26 974
rect 26 1008 92 1024
rect 26 974 42 1008
rect 76 974 92 1008
rect 26 958 92 974
rect 144 1008 210 1024
rect 144 974 160 1008
rect 194 974 210 1008
rect 144 958 210 974
rect 262 1008 328 1024
rect 262 974 278 1008
rect 312 974 328 1008
rect 262 958 328 974
rect 380 1008 446 1024
rect 380 974 396 1008
rect 430 974 446 1008
rect 380 958 446 974
rect 498 1008 564 1024
rect 498 974 514 1008
rect 548 974 564 1008
rect 498 958 564 974
rect -561 936 -501 958
rect -443 936 -383 958
rect -325 936 -265 958
rect -207 936 -147 958
rect -89 936 -29 958
rect 29 936 89 958
rect 147 936 207 958
rect 265 936 325 958
rect 383 936 443 958
rect 501 936 561 958
rect -561 714 -501 736
rect -443 714 -383 736
rect -325 714 -265 736
rect -207 714 -147 736
rect -89 714 -29 736
rect 29 714 89 736
rect 147 714 207 736
rect 265 714 325 736
rect 383 714 443 736
rect 501 714 561 736
rect -564 698 -498 714
rect -564 664 -548 698
rect -514 664 -498 698
rect -564 648 -498 664
rect -446 698 -380 714
rect -446 664 -430 698
rect -396 664 -380 698
rect -446 648 -380 664
rect -328 698 -262 714
rect -328 664 -312 698
rect -278 664 -262 698
rect -328 648 -262 664
rect -210 698 -144 714
rect -210 664 -194 698
rect -160 664 -144 698
rect -210 648 -144 664
rect -92 698 -26 714
rect -92 664 -76 698
rect -42 664 -26 698
rect -92 648 -26 664
rect 26 698 92 714
rect 26 664 42 698
rect 76 664 92 698
rect 26 648 92 664
rect 144 698 210 714
rect 144 664 160 698
rect 194 664 210 698
rect 144 648 210 664
rect 262 698 328 714
rect 262 664 278 698
rect 312 664 328 698
rect 262 648 328 664
rect 380 698 446 714
rect 380 664 396 698
rect 430 664 446 698
rect 380 648 446 664
rect 498 698 564 714
rect 498 664 514 698
rect 548 664 564 698
rect 498 648 564 664
rect -564 590 -498 606
rect -564 556 -548 590
rect -514 556 -498 590
rect -564 540 -498 556
rect -446 590 -380 606
rect -446 556 -430 590
rect -396 556 -380 590
rect -446 540 -380 556
rect -328 590 -262 606
rect -328 556 -312 590
rect -278 556 -262 590
rect -328 540 -262 556
rect -210 590 -144 606
rect -210 556 -194 590
rect -160 556 -144 590
rect -210 540 -144 556
rect -92 590 -26 606
rect -92 556 -76 590
rect -42 556 -26 590
rect -92 540 -26 556
rect 26 590 92 606
rect 26 556 42 590
rect 76 556 92 590
rect 26 540 92 556
rect 144 590 210 606
rect 144 556 160 590
rect 194 556 210 590
rect 144 540 210 556
rect 262 590 328 606
rect 262 556 278 590
rect 312 556 328 590
rect 262 540 328 556
rect 380 590 446 606
rect 380 556 396 590
rect 430 556 446 590
rect 380 540 446 556
rect 498 590 564 606
rect 498 556 514 590
rect 548 556 564 590
rect 498 540 564 556
rect -561 518 -501 540
rect -443 518 -383 540
rect -325 518 -265 540
rect -207 518 -147 540
rect -89 518 -29 540
rect 29 518 89 540
rect 147 518 207 540
rect 265 518 325 540
rect 383 518 443 540
rect 501 518 561 540
rect -561 296 -501 318
rect -443 296 -383 318
rect -325 296 -265 318
rect -207 296 -147 318
rect -89 296 -29 318
rect 29 296 89 318
rect 147 296 207 318
rect 265 296 325 318
rect 383 296 443 318
rect 501 296 561 318
rect -564 280 -498 296
rect -564 246 -548 280
rect -514 246 -498 280
rect -564 230 -498 246
rect -446 280 -380 296
rect -446 246 -430 280
rect -396 246 -380 280
rect -446 230 -380 246
rect -328 280 -262 296
rect -328 246 -312 280
rect -278 246 -262 280
rect -328 230 -262 246
rect -210 280 -144 296
rect -210 246 -194 280
rect -160 246 -144 280
rect -210 230 -144 246
rect -92 280 -26 296
rect -92 246 -76 280
rect -42 246 -26 280
rect -92 230 -26 246
rect 26 280 92 296
rect 26 246 42 280
rect 76 246 92 280
rect 26 230 92 246
rect 144 280 210 296
rect 144 246 160 280
rect 194 246 210 280
rect 144 230 210 246
rect 262 280 328 296
rect 262 246 278 280
rect 312 246 328 280
rect 262 230 328 246
rect 380 280 446 296
rect 380 246 396 280
rect 430 246 446 280
rect 380 230 446 246
rect 498 280 564 296
rect 498 246 514 280
rect 548 246 564 280
rect 498 230 564 246
rect -564 172 -498 188
rect -564 138 -548 172
rect -514 138 -498 172
rect -564 122 -498 138
rect -446 172 -380 188
rect -446 138 -430 172
rect -396 138 -380 172
rect -446 122 -380 138
rect -328 172 -262 188
rect -328 138 -312 172
rect -278 138 -262 172
rect -328 122 -262 138
rect -210 172 -144 188
rect -210 138 -194 172
rect -160 138 -144 172
rect -210 122 -144 138
rect -92 172 -26 188
rect -92 138 -76 172
rect -42 138 -26 172
rect -92 122 -26 138
rect 26 172 92 188
rect 26 138 42 172
rect 76 138 92 172
rect 26 122 92 138
rect 144 172 210 188
rect 144 138 160 172
rect 194 138 210 172
rect 144 122 210 138
rect 262 172 328 188
rect 262 138 278 172
rect 312 138 328 172
rect 262 122 328 138
rect 380 172 446 188
rect 380 138 396 172
rect 430 138 446 172
rect 380 122 446 138
rect 498 172 564 188
rect 498 138 514 172
rect 548 138 564 172
rect 498 122 564 138
rect -561 100 -501 122
rect -443 100 -383 122
rect -325 100 -265 122
rect -207 100 -147 122
rect -89 100 -29 122
rect 29 100 89 122
rect 147 100 207 122
rect 265 100 325 122
rect 383 100 443 122
rect 501 100 561 122
rect -561 -122 -501 -100
rect -443 -122 -383 -100
rect -325 -122 -265 -100
rect -207 -122 -147 -100
rect -89 -122 -29 -100
rect 29 -122 89 -100
rect 147 -122 207 -100
rect 265 -122 325 -100
rect 383 -122 443 -100
rect 501 -122 561 -100
rect -564 -138 -498 -122
rect -564 -172 -548 -138
rect -514 -172 -498 -138
rect -564 -188 -498 -172
rect -446 -138 -380 -122
rect -446 -172 -430 -138
rect -396 -172 -380 -138
rect -446 -188 -380 -172
rect -328 -138 -262 -122
rect -328 -172 -312 -138
rect -278 -172 -262 -138
rect -328 -188 -262 -172
rect -210 -138 -144 -122
rect -210 -172 -194 -138
rect -160 -172 -144 -138
rect -210 -188 -144 -172
rect -92 -138 -26 -122
rect -92 -172 -76 -138
rect -42 -172 -26 -138
rect -92 -188 -26 -172
rect 26 -138 92 -122
rect 26 -172 42 -138
rect 76 -172 92 -138
rect 26 -188 92 -172
rect 144 -138 210 -122
rect 144 -172 160 -138
rect 194 -172 210 -138
rect 144 -188 210 -172
rect 262 -138 328 -122
rect 262 -172 278 -138
rect 312 -172 328 -138
rect 262 -188 328 -172
rect 380 -138 446 -122
rect 380 -172 396 -138
rect 430 -172 446 -138
rect 380 -188 446 -172
rect 498 -138 564 -122
rect 498 -172 514 -138
rect 548 -172 564 -138
rect 498 -188 564 -172
rect -564 -246 -498 -230
rect -564 -280 -548 -246
rect -514 -280 -498 -246
rect -564 -296 -498 -280
rect -446 -246 -380 -230
rect -446 -280 -430 -246
rect -396 -280 -380 -246
rect -446 -296 -380 -280
rect -328 -246 -262 -230
rect -328 -280 -312 -246
rect -278 -280 -262 -246
rect -328 -296 -262 -280
rect -210 -246 -144 -230
rect -210 -280 -194 -246
rect -160 -280 -144 -246
rect -210 -296 -144 -280
rect -92 -246 -26 -230
rect -92 -280 -76 -246
rect -42 -280 -26 -246
rect -92 -296 -26 -280
rect 26 -246 92 -230
rect 26 -280 42 -246
rect 76 -280 92 -246
rect 26 -296 92 -280
rect 144 -246 210 -230
rect 144 -280 160 -246
rect 194 -280 210 -246
rect 144 -296 210 -280
rect 262 -246 328 -230
rect 262 -280 278 -246
rect 312 -280 328 -246
rect 262 -296 328 -280
rect 380 -246 446 -230
rect 380 -280 396 -246
rect 430 -280 446 -246
rect 380 -296 446 -280
rect 498 -246 564 -230
rect 498 -280 514 -246
rect 548 -280 564 -246
rect 498 -296 564 -280
rect -561 -318 -501 -296
rect -443 -318 -383 -296
rect -325 -318 -265 -296
rect -207 -318 -147 -296
rect -89 -318 -29 -296
rect 29 -318 89 -296
rect 147 -318 207 -296
rect 265 -318 325 -296
rect 383 -318 443 -296
rect 501 -318 561 -296
rect -561 -540 -501 -518
rect -443 -540 -383 -518
rect -325 -540 -265 -518
rect -207 -540 -147 -518
rect -89 -540 -29 -518
rect 29 -540 89 -518
rect 147 -540 207 -518
rect 265 -540 325 -518
rect 383 -540 443 -518
rect 501 -540 561 -518
rect -564 -556 -498 -540
rect -564 -590 -548 -556
rect -514 -590 -498 -556
rect -564 -606 -498 -590
rect -446 -556 -380 -540
rect -446 -590 -430 -556
rect -396 -590 -380 -556
rect -446 -606 -380 -590
rect -328 -556 -262 -540
rect -328 -590 -312 -556
rect -278 -590 -262 -556
rect -328 -606 -262 -590
rect -210 -556 -144 -540
rect -210 -590 -194 -556
rect -160 -590 -144 -556
rect -210 -606 -144 -590
rect -92 -556 -26 -540
rect -92 -590 -76 -556
rect -42 -590 -26 -556
rect -92 -606 -26 -590
rect 26 -556 92 -540
rect 26 -590 42 -556
rect 76 -590 92 -556
rect 26 -606 92 -590
rect 144 -556 210 -540
rect 144 -590 160 -556
rect 194 -590 210 -556
rect 144 -606 210 -590
rect 262 -556 328 -540
rect 262 -590 278 -556
rect 312 -590 328 -556
rect 262 -606 328 -590
rect 380 -556 446 -540
rect 380 -590 396 -556
rect 430 -590 446 -556
rect 380 -606 446 -590
rect 498 -556 564 -540
rect 498 -590 514 -556
rect 548 -590 564 -556
rect 498 -606 564 -590
rect -564 -664 -498 -648
rect -564 -698 -548 -664
rect -514 -698 -498 -664
rect -564 -714 -498 -698
rect -446 -664 -380 -648
rect -446 -698 -430 -664
rect -396 -698 -380 -664
rect -446 -714 -380 -698
rect -328 -664 -262 -648
rect -328 -698 -312 -664
rect -278 -698 -262 -664
rect -328 -714 -262 -698
rect -210 -664 -144 -648
rect -210 -698 -194 -664
rect -160 -698 -144 -664
rect -210 -714 -144 -698
rect -92 -664 -26 -648
rect -92 -698 -76 -664
rect -42 -698 -26 -664
rect -92 -714 -26 -698
rect 26 -664 92 -648
rect 26 -698 42 -664
rect 76 -698 92 -664
rect 26 -714 92 -698
rect 144 -664 210 -648
rect 144 -698 160 -664
rect 194 -698 210 -664
rect 144 -714 210 -698
rect 262 -664 328 -648
rect 262 -698 278 -664
rect 312 -698 328 -664
rect 262 -714 328 -698
rect 380 -664 446 -648
rect 380 -698 396 -664
rect 430 -698 446 -664
rect 380 -714 446 -698
rect 498 -664 564 -648
rect 498 -698 514 -664
rect 548 -698 564 -664
rect 498 -714 564 -698
rect -561 -736 -501 -714
rect -443 -736 -383 -714
rect -325 -736 -265 -714
rect -207 -736 -147 -714
rect -89 -736 -29 -714
rect 29 -736 89 -714
rect 147 -736 207 -714
rect 265 -736 325 -714
rect 383 -736 443 -714
rect 501 -736 561 -714
rect -561 -958 -501 -936
rect -443 -958 -383 -936
rect -325 -958 -265 -936
rect -207 -958 -147 -936
rect -89 -958 -29 -936
rect 29 -958 89 -936
rect 147 -958 207 -936
rect 265 -958 325 -936
rect 383 -958 443 -936
rect 501 -958 561 -936
rect -564 -974 -498 -958
rect -564 -1008 -548 -974
rect -514 -1008 -498 -974
rect -564 -1024 -498 -1008
rect -446 -974 -380 -958
rect -446 -1008 -430 -974
rect -396 -1008 -380 -974
rect -446 -1024 -380 -1008
rect -328 -974 -262 -958
rect -328 -1008 -312 -974
rect -278 -1008 -262 -974
rect -328 -1024 -262 -1008
rect -210 -974 -144 -958
rect -210 -1008 -194 -974
rect -160 -1008 -144 -974
rect -210 -1024 -144 -1008
rect -92 -974 -26 -958
rect -92 -1008 -76 -974
rect -42 -1008 -26 -974
rect -92 -1024 -26 -1008
rect 26 -974 92 -958
rect 26 -1008 42 -974
rect 76 -1008 92 -974
rect 26 -1024 92 -1008
rect 144 -974 210 -958
rect 144 -1008 160 -974
rect 194 -1008 210 -974
rect 144 -1024 210 -1008
rect 262 -974 328 -958
rect 262 -1008 278 -974
rect 312 -1008 328 -974
rect 262 -1024 328 -1008
rect 380 -974 446 -958
rect 380 -1008 396 -974
rect 430 -1008 446 -974
rect 380 -1024 446 -1008
rect 498 -974 564 -958
rect 498 -1008 514 -974
rect 548 -1008 564 -974
rect 498 -1024 564 -1008
<< polycont >>
rect -548 974 -514 1008
rect -430 974 -396 1008
rect -312 974 -278 1008
rect -194 974 -160 1008
rect -76 974 -42 1008
rect 42 974 76 1008
rect 160 974 194 1008
rect 278 974 312 1008
rect 396 974 430 1008
rect 514 974 548 1008
rect -548 664 -514 698
rect -430 664 -396 698
rect -312 664 -278 698
rect -194 664 -160 698
rect -76 664 -42 698
rect 42 664 76 698
rect 160 664 194 698
rect 278 664 312 698
rect 396 664 430 698
rect 514 664 548 698
rect -548 556 -514 590
rect -430 556 -396 590
rect -312 556 -278 590
rect -194 556 -160 590
rect -76 556 -42 590
rect 42 556 76 590
rect 160 556 194 590
rect 278 556 312 590
rect 396 556 430 590
rect 514 556 548 590
rect -548 246 -514 280
rect -430 246 -396 280
rect -312 246 -278 280
rect -194 246 -160 280
rect -76 246 -42 280
rect 42 246 76 280
rect 160 246 194 280
rect 278 246 312 280
rect 396 246 430 280
rect 514 246 548 280
rect -548 138 -514 172
rect -430 138 -396 172
rect -312 138 -278 172
rect -194 138 -160 172
rect -76 138 -42 172
rect 42 138 76 172
rect 160 138 194 172
rect 278 138 312 172
rect 396 138 430 172
rect 514 138 548 172
rect -548 -172 -514 -138
rect -430 -172 -396 -138
rect -312 -172 -278 -138
rect -194 -172 -160 -138
rect -76 -172 -42 -138
rect 42 -172 76 -138
rect 160 -172 194 -138
rect 278 -172 312 -138
rect 396 -172 430 -138
rect 514 -172 548 -138
rect -548 -280 -514 -246
rect -430 -280 -396 -246
rect -312 -280 -278 -246
rect -194 -280 -160 -246
rect -76 -280 -42 -246
rect 42 -280 76 -246
rect 160 -280 194 -246
rect 278 -280 312 -246
rect 396 -280 430 -246
rect 514 -280 548 -246
rect -548 -590 -514 -556
rect -430 -590 -396 -556
rect -312 -590 -278 -556
rect -194 -590 -160 -556
rect -76 -590 -42 -556
rect 42 -590 76 -556
rect 160 -590 194 -556
rect 278 -590 312 -556
rect 396 -590 430 -556
rect 514 -590 548 -556
rect -548 -698 -514 -664
rect -430 -698 -396 -664
rect -312 -698 -278 -664
rect -194 -698 -160 -664
rect -76 -698 -42 -664
rect 42 -698 76 -664
rect 160 -698 194 -664
rect 278 -698 312 -664
rect 396 -698 430 -664
rect 514 -698 548 -664
rect -548 -1008 -514 -974
rect -430 -1008 -396 -974
rect -312 -1008 -278 -974
rect -194 -1008 -160 -974
rect -76 -1008 -42 -974
rect 42 -1008 76 -974
rect 160 -1008 194 -974
rect 278 -1008 312 -974
rect 396 -1008 430 -974
rect 514 -1008 548 -974
<< locali >>
rect -721 1076 -625 1110
rect 625 1076 721 1110
rect -721 1014 -687 1076
rect 687 1014 721 1076
rect -564 974 -548 1008
rect -514 974 -498 1008
rect -446 974 -430 1008
rect -396 974 -380 1008
rect -328 974 -312 1008
rect -278 974 -262 1008
rect -210 974 -194 1008
rect -160 974 -144 1008
rect -92 974 -76 1008
rect -42 974 -26 1008
rect 26 974 42 1008
rect 76 974 92 1008
rect 144 974 160 1008
rect 194 974 210 1008
rect 262 974 278 1008
rect 312 974 328 1008
rect 380 974 396 1008
rect 430 974 446 1008
rect 498 974 514 1008
rect 548 974 564 1008
rect -607 924 -573 940
rect -607 732 -573 748
rect -489 924 -455 940
rect -489 732 -455 748
rect -371 924 -337 940
rect -371 732 -337 748
rect -253 924 -219 940
rect -253 732 -219 748
rect -135 924 -101 940
rect -135 732 -101 748
rect -17 924 17 940
rect -17 732 17 748
rect 101 924 135 940
rect 101 732 135 748
rect 219 924 253 940
rect 219 732 253 748
rect 337 924 371 940
rect 337 732 371 748
rect 455 924 489 940
rect 455 732 489 748
rect 573 924 607 940
rect 573 732 607 748
rect -564 664 -548 698
rect -514 664 -498 698
rect -446 664 -430 698
rect -396 664 -380 698
rect -328 664 -312 698
rect -278 664 -262 698
rect -210 664 -194 698
rect -160 664 -144 698
rect -92 664 -76 698
rect -42 664 -26 698
rect 26 664 42 698
rect 76 664 92 698
rect 144 664 160 698
rect 194 664 210 698
rect 262 664 278 698
rect 312 664 328 698
rect 380 664 396 698
rect 430 664 446 698
rect 498 664 514 698
rect 548 664 564 698
rect -564 556 -548 590
rect -514 556 -498 590
rect -446 556 -430 590
rect -396 556 -380 590
rect -328 556 -312 590
rect -278 556 -262 590
rect -210 556 -194 590
rect -160 556 -144 590
rect -92 556 -76 590
rect -42 556 -26 590
rect 26 556 42 590
rect 76 556 92 590
rect 144 556 160 590
rect 194 556 210 590
rect 262 556 278 590
rect 312 556 328 590
rect 380 556 396 590
rect 430 556 446 590
rect 498 556 514 590
rect 548 556 564 590
rect -607 506 -573 522
rect -607 314 -573 330
rect -489 506 -455 522
rect -489 314 -455 330
rect -371 506 -337 522
rect -371 314 -337 330
rect -253 506 -219 522
rect -253 314 -219 330
rect -135 506 -101 522
rect -135 314 -101 330
rect -17 506 17 522
rect -17 314 17 330
rect 101 506 135 522
rect 101 314 135 330
rect 219 506 253 522
rect 219 314 253 330
rect 337 506 371 522
rect 337 314 371 330
rect 455 506 489 522
rect 455 314 489 330
rect 573 506 607 522
rect 573 314 607 330
rect -564 246 -548 280
rect -514 246 -498 280
rect -446 246 -430 280
rect -396 246 -380 280
rect -328 246 -312 280
rect -278 246 -262 280
rect -210 246 -194 280
rect -160 246 -144 280
rect -92 246 -76 280
rect -42 246 -26 280
rect 26 246 42 280
rect 76 246 92 280
rect 144 246 160 280
rect 194 246 210 280
rect 262 246 278 280
rect 312 246 328 280
rect 380 246 396 280
rect 430 246 446 280
rect 498 246 514 280
rect 548 246 564 280
rect -564 138 -548 172
rect -514 138 -498 172
rect -446 138 -430 172
rect -396 138 -380 172
rect -328 138 -312 172
rect -278 138 -262 172
rect -210 138 -194 172
rect -160 138 -144 172
rect -92 138 -76 172
rect -42 138 -26 172
rect 26 138 42 172
rect 76 138 92 172
rect 144 138 160 172
rect 194 138 210 172
rect 262 138 278 172
rect 312 138 328 172
rect 380 138 396 172
rect 430 138 446 172
rect 498 138 514 172
rect 548 138 564 172
rect -607 88 -573 104
rect -607 -104 -573 -88
rect -489 88 -455 104
rect -489 -104 -455 -88
rect -371 88 -337 104
rect -371 -104 -337 -88
rect -253 88 -219 104
rect -253 -104 -219 -88
rect -135 88 -101 104
rect -135 -104 -101 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 101 88 135 104
rect 101 -104 135 -88
rect 219 88 253 104
rect 219 -104 253 -88
rect 337 88 371 104
rect 337 -104 371 -88
rect 455 88 489 104
rect 455 -104 489 -88
rect 573 88 607 104
rect 573 -104 607 -88
rect -564 -172 -548 -138
rect -514 -172 -498 -138
rect -446 -172 -430 -138
rect -396 -172 -380 -138
rect -328 -172 -312 -138
rect -278 -172 -262 -138
rect -210 -172 -194 -138
rect -160 -172 -144 -138
rect -92 -172 -76 -138
rect -42 -172 -26 -138
rect 26 -172 42 -138
rect 76 -172 92 -138
rect 144 -172 160 -138
rect 194 -172 210 -138
rect 262 -172 278 -138
rect 312 -172 328 -138
rect 380 -172 396 -138
rect 430 -172 446 -138
rect 498 -172 514 -138
rect 548 -172 564 -138
rect -564 -280 -548 -246
rect -514 -280 -498 -246
rect -446 -280 -430 -246
rect -396 -280 -380 -246
rect -328 -280 -312 -246
rect -278 -280 -262 -246
rect -210 -280 -194 -246
rect -160 -280 -144 -246
rect -92 -280 -76 -246
rect -42 -280 -26 -246
rect 26 -280 42 -246
rect 76 -280 92 -246
rect 144 -280 160 -246
rect 194 -280 210 -246
rect 262 -280 278 -246
rect 312 -280 328 -246
rect 380 -280 396 -246
rect 430 -280 446 -246
rect 498 -280 514 -246
rect 548 -280 564 -246
rect -607 -330 -573 -314
rect -607 -522 -573 -506
rect -489 -330 -455 -314
rect -489 -522 -455 -506
rect -371 -330 -337 -314
rect -371 -522 -337 -506
rect -253 -330 -219 -314
rect -253 -522 -219 -506
rect -135 -330 -101 -314
rect -135 -522 -101 -506
rect -17 -330 17 -314
rect -17 -522 17 -506
rect 101 -330 135 -314
rect 101 -522 135 -506
rect 219 -330 253 -314
rect 219 -522 253 -506
rect 337 -330 371 -314
rect 337 -522 371 -506
rect 455 -330 489 -314
rect 455 -522 489 -506
rect 573 -330 607 -314
rect 573 -522 607 -506
rect -564 -590 -548 -556
rect -514 -590 -498 -556
rect -446 -590 -430 -556
rect -396 -590 -380 -556
rect -328 -590 -312 -556
rect -278 -590 -262 -556
rect -210 -590 -194 -556
rect -160 -590 -144 -556
rect -92 -590 -76 -556
rect -42 -590 -26 -556
rect 26 -590 42 -556
rect 76 -590 92 -556
rect 144 -590 160 -556
rect 194 -590 210 -556
rect 262 -590 278 -556
rect 312 -590 328 -556
rect 380 -590 396 -556
rect 430 -590 446 -556
rect 498 -590 514 -556
rect 548 -590 564 -556
rect -564 -698 -548 -664
rect -514 -698 -498 -664
rect -446 -698 -430 -664
rect -396 -698 -380 -664
rect -328 -698 -312 -664
rect -278 -698 -262 -664
rect -210 -698 -194 -664
rect -160 -698 -144 -664
rect -92 -698 -76 -664
rect -42 -698 -26 -664
rect 26 -698 42 -664
rect 76 -698 92 -664
rect 144 -698 160 -664
rect 194 -698 210 -664
rect 262 -698 278 -664
rect 312 -698 328 -664
rect 380 -698 396 -664
rect 430 -698 446 -664
rect 498 -698 514 -664
rect 548 -698 564 -664
rect -607 -748 -573 -732
rect -607 -940 -573 -924
rect -489 -748 -455 -732
rect -489 -940 -455 -924
rect -371 -748 -337 -732
rect -371 -940 -337 -924
rect -253 -748 -219 -732
rect -253 -940 -219 -924
rect -135 -748 -101 -732
rect -135 -940 -101 -924
rect -17 -748 17 -732
rect -17 -940 17 -924
rect 101 -748 135 -732
rect 101 -940 135 -924
rect 219 -748 253 -732
rect 219 -940 253 -924
rect 337 -748 371 -732
rect 337 -940 371 -924
rect 455 -748 489 -732
rect 455 -940 489 -924
rect 573 -748 607 -732
rect 573 -940 607 -924
rect -564 -1008 -548 -974
rect -514 -1008 -498 -974
rect -446 -1008 -430 -974
rect -396 -1008 -380 -974
rect -328 -1008 -312 -974
rect -278 -1008 -262 -974
rect -210 -1008 -194 -974
rect -160 -1008 -144 -974
rect -92 -1008 -76 -974
rect -42 -1008 -26 -974
rect 26 -1008 42 -974
rect 76 -1008 92 -974
rect 144 -1008 160 -974
rect 194 -1008 210 -974
rect 262 -1008 278 -974
rect 312 -1008 328 -974
rect 380 -1008 396 -974
rect 430 -1008 446 -974
rect 498 -1008 514 -974
rect 548 -1008 564 -974
rect -721 -1076 -687 -1014
rect 687 -1076 721 -1014
rect -721 -1110 -625 -1076
rect 625 -1110 721 -1076
<< viali >>
rect -548 974 -514 1008
rect -430 974 -396 1008
rect -312 974 -278 1008
rect -194 974 -160 1008
rect -76 974 -42 1008
rect 42 974 76 1008
rect 160 974 194 1008
rect 278 974 312 1008
rect 396 974 430 1008
rect 514 974 548 1008
rect -607 748 -573 924
rect -489 748 -455 924
rect -371 748 -337 924
rect -253 748 -219 924
rect -135 748 -101 924
rect -17 748 17 924
rect 101 748 135 924
rect 219 748 253 924
rect 337 748 371 924
rect 455 748 489 924
rect 573 748 607 924
rect -548 664 -514 698
rect -430 664 -396 698
rect -312 664 -278 698
rect -194 664 -160 698
rect -76 664 -42 698
rect 42 664 76 698
rect 160 664 194 698
rect 278 664 312 698
rect 396 664 430 698
rect 514 664 548 698
rect -548 556 -514 590
rect -430 556 -396 590
rect -312 556 -278 590
rect -194 556 -160 590
rect -76 556 -42 590
rect 42 556 76 590
rect 160 556 194 590
rect 278 556 312 590
rect 396 556 430 590
rect 514 556 548 590
rect -607 330 -573 506
rect -489 330 -455 506
rect -371 330 -337 506
rect -253 330 -219 506
rect -135 330 -101 506
rect -17 330 17 506
rect 101 330 135 506
rect 219 330 253 506
rect 337 330 371 506
rect 455 330 489 506
rect 573 330 607 506
rect -548 246 -514 280
rect -430 246 -396 280
rect -312 246 -278 280
rect -194 246 -160 280
rect -76 246 -42 280
rect 42 246 76 280
rect 160 246 194 280
rect 278 246 312 280
rect 396 246 430 280
rect 514 246 548 280
rect -548 138 -514 172
rect -430 138 -396 172
rect -312 138 -278 172
rect -194 138 -160 172
rect -76 138 -42 172
rect 42 138 76 172
rect 160 138 194 172
rect 278 138 312 172
rect 396 138 430 172
rect 514 138 548 172
rect -607 -88 -573 88
rect -489 -88 -455 88
rect -371 -88 -337 88
rect -253 -88 -219 88
rect -135 -88 -101 88
rect -17 -88 17 88
rect 101 -88 135 88
rect 219 -88 253 88
rect 337 -88 371 88
rect 455 -88 489 88
rect 573 -88 607 88
rect -548 -172 -514 -138
rect -430 -172 -396 -138
rect -312 -172 -278 -138
rect -194 -172 -160 -138
rect -76 -172 -42 -138
rect 42 -172 76 -138
rect 160 -172 194 -138
rect 278 -172 312 -138
rect 396 -172 430 -138
rect 514 -172 548 -138
rect -548 -280 -514 -246
rect -430 -280 -396 -246
rect -312 -280 -278 -246
rect -194 -280 -160 -246
rect -76 -280 -42 -246
rect 42 -280 76 -246
rect 160 -280 194 -246
rect 278 -280 312 -246
rect 396 -280 430 -246
rect 514 -280 548 -246
rect -607 -506 -573 -330
rect -489 -506 -455 -330
rect -371 -506 -337 -330
rect -253 -506 -219 -330
rect -135 -506 -101 -330
rect -17 -506 17 -330
rect 101 -506 135 -330
rect 219 -506 253 -330
rect 337 -506 371 -330
rect 455 -506 489 -330
rect 573 -506 607 -330
rect -548 -590 -514 -556
rect -430 -590 -396 -556
rect -312 -590 -278 -556
rect -194 -590 -160 -556
rect -76 -590 -42 -556
rect 42 -590 76 -556
rect 160 -590 194 -556
rect 278 -590 312 -556
rect 396 -590 430 -556
rect 514 -590 548 -556
rect -548 -698 -514 -664
rect -430 -698 -396 -664
rect -312 -698 -278 -664
rect -194 -698 -160 -664
rect -76 -698 -42 -664
rect 42 -698 76 -664
rect 160 -698 194 -664
rect 278 -698 312 -664
rect 396 -698 430 -664
rect 514 -698 548 -664
rect -607 -924 -573 -748
rect -489 -924 -455 -748
rect -371 -924 -337 -748
rect -253 -924 -219 -748
rect -135 -924 -101 -748
rect -17 -924 17 -748
rect 101 -924 135 -748
rect 219 -924 253 -748
rect 337 -924 371 -748
rect 455 -924 489 -748
rect 573 -924 607 -748
rect -548 -1008 -514 -974
rect -430 -1008 -396 -974
rect -312 -1008 -278 -974
rect -194 -1008 -160 -974
rect -76 -1008 -42 -974
rect 42 -1008 76 -974
rect 160 -1008 194 -974
rect 278 -1008 312 -974
rect 396 -1008 430 -974
rect 514 -1008 548 -974
<< metal1 >>
rect -560 1008 -502 1014
rect -560 974 -548 1008
rect -514 974 -502 1008
rect -560 968 -502 974
rect -442 1008 -384 1014
rect -442 974 -430 1008
rect -396 974 -384 1008
rect -442 968 -384 974
rect -324 1008 -266 1014
rect -324 974 -312 1008
rect -278 974 -266 1008
rect -324 968 -266 974
rect -206 1008 -148 1014
rect -206 974 -194 1008
rect -160 974 -148 1008
rect -206 968 -148 974
rect -88 1008 -30 1014
rect -88 974 -76 1008
rect -42 974 -30 1008
rect -88 968 -30 974
rect 30 1008 88 1014
rect 30 974 42 1008
rect 76 974 88 1008
rect 30 968 88 974
rect 148 1008 206 1014
rect 148 974 160 1008
rect 194 974 206 1008
rect 148 968 206 974
rect 266 1008 324 1014
rect 266 974 278 1008
rect 312 974 324 1008
rect 266 968 324 974
rect 384 1008 442 1014
rect 384 974 396 1008
rect 430 974 442 1008
rect 384 968 442 974
rect 502 1008 560 1014
rect 502 974 514 1008
rect 548 974 560 1008
rect 502 968 560 974
rect -613 924 -567 936
rect -613 748 -607 924
rect -573 748 -567 924
rect -613 736 -567 748
rect -495 924 -449 936
rect -495 748 -489 924
rect -455 748 -449 924
rect -495 736 -449 748
rect -377 924 -331 936
rect -377 748 -371 924
rect -337 748 -331 924
rect -377 736 -331 748
rect -259 924 -213 936
rect -259 748 -253 924
rect -219 748 -213 924
rect -259 736 -213 748
rect -141 924 -95 936
rect -141 748 -135 924
rect -101 748 -95 924
rect -141 736 -95 748
rect -23 924 23 936
rect -23 748 -17 924
rect 17 748 23 924
rect -23 736 23 748
rect 95 924 141 936
rect 95 748 101 924
rect 135 748 141 924
rect 95 736 141 748
rect 213 924 259 936
rect 213 748 219 924
rect 253 748 259 924
rect 213 736 259 748
rect 331 924 377 936
rect 331 748 337 924
rect 371 748 377 924
rect 331 736 377 748
rect 449 924 495 936
rect 449 748 455 924
rect 489 748 495 924
rect 449 736 495 748
rect 567 924 613 936
rect 567 748 573 924
rect 607 748 613 924
rect 567 736 613 748
rect -560 698 -502 704
rect -560 664 -548 698
rect -514 664 -502 698
rect -560 658 -502 664
rect -442 698 -384 704
rect -442 664 -430 698
rect -396 664 -384 698
rect -442 658 -384 664
rect -324 698 -266 704
rect -324 664 -312 698
rect -278 664 -266 698
rect -324 658 -266 664
rect -206 698 -148 704
rect -206 664 -194 698
rect -160 664 -148 698
rect -206 658 -148 664
rect -88 698 -30 704
rect -88 664 -76 698
rect -42 664 -30 698
rect -88 658 -30 664
rect 30 698 88 704
rect 30 664 42 698
rect 76 664 88 698
rect 30 658 88 664
rect 148 698 206 704
rect 148 664 160 698
rect 194 664 206 698
rect 148 658 206 664
rect 266 698 324 704
rect 266 664 278 698
rect 312 664 324 698
rect 266 658 324 664
rect 384 698 442 704
rect 384 664 396 698
rect 430 664 442 698
rect 384 658 442 664
rect 502 698 560 704
rect 502 664 514 698
rect 548 664 560 698
rect 502 658 560 664
rect -560 590 -502 596
rect -560 556 -548 590
rect -514 556 -502 590
rect -560 550 -502 556
rect -442 590 -384 596
rect -442 556 -430 590
rect -396 556 -384 590
rect -442 550 -384 556
rect -324 590 -266 596
rect -324 556 -312 590
rect -278 556 -266 590
rect -324 550 -266 556
rect -206 590 -148 596
rect -206 556 -194 590
rect -160 556 -148 590
rect -206 550 -148 556
rect -88 590 -30 596
rect -88 556 -76 590
rect -42 556 -30 590
rect -88 550 -30 556
rect 30 590 88 596
rect 30 556 42 590
rect 76 556 88 590
rect 30 550 88 556
rect 148 590 206 596
rect 148 556 160 590
rect 194 556 206 590
rect 148 550 206 556
rect 266 590 324 596
rect 266 556 278 590
rect 312 556 324 590
rect 266 550 324 556
rect 384 590 442 596
rect 384 556 396 590
rect 430 556 442 590
rect 384 550 442 556
rect 502 590 560 596
rect 502 556 514 590
rect 548 556 560 590
rect 502 550 560 556
rect -613 506 -567 518
rect -613 330 -607 506
rect -573 330 -567 506
rect -613 318 -567 330
rect -495 506 -449 518
rect -495 330 -489 506
rect -455 330 -449 506
rect -495 318 -449 330
rect -377 506 -331 518
rect -377 330 -371 506
rect -337 330 -331 506
rect -377 318 -331 330
rect -259 506 -213 518
rect -259 330 -253 506
rect -219 330 -213 506
rect -259 318 -213 330
rect -141 506 -95 518
rect -141 330 -135 506
rect -101 330 -95 506
rect -141 318 -95 330
rect -23 506 23 518
rect -23 330 -17 506
rect 17 330 23 506
rect -23 318 23 330
rect 95 506 141 518
rect 95 330 101 506
rect 135 330 141 506
rect 95 318 141 330
rect 213 506 259 518
rect 213 330 219 506
rect 253 330 259 506
rect 213 318 259 330
rect 331 506 377 518
rect 331 330 337 506
rect 371 330 377 506
rect 331 318 377 330
rect 449 506 495 518
rect 449 330 455 506
rect 489 330 495 506
rect 449 318 495 330
rect 567 506 613 518
rect 567 330 573 506
rect 607 330 613 506
rect 567 318 613 330
rect -560 280 -502 286
rect -560 246 -548 280
rect -514 246 -502 280
rect -560 240 -502 246
rect -442 280 -384 286
rect -442 246 -430 280
rect -396 246 -384 280
rect -442 240 -384 246
rect -324 280 -266 286
rect -324 246 -312 280
rect -278 246 -266 280
rect -324 240 -266 246
rect -206 280 -148 286
rect -206 246 -194 280
rect -160 246 -148 280
rect -206 240 -148 246
rect -88 280 -30 286
rect -88 246 -76 280
rect -42 246 -30 280
rect -88 240 -30 246
rect 30 280 88 286
rect 30 246 42 280
rect 76 246 88 280
rect 30 240 88 246
rect 148 280 206 286
rect 148 246 160 280
rect 194 246 206 280
rect 148 240 206 246
rect 266 280 324 286
rect 266 246 278 280
rect 312 246 324 280
rect 266 240 324 246
rect 384 280 442 286
rect 384 246 396 280
rect 430 246 442 280
rect 384 240 442 246
rect 502 280 560 286
rect 502 246 514 280
rect 548 246 560 280
rect 502 240 560 246
rect -560 172 -502 178
rect -560 138 -548 172
rect -514 138 -502 172
rect -560 132 -502 138
rect -442 172 -384 178
rect -442 138 -430 172
rect -396 138 -384 172
rect -442 132 -384 138
rect -324 172 -266 178
rect -324 138 -312 172
rect -278 138 -266 172
rect -324 132 -266 138
rect -206 172 -148 178
rect -206 138 -194 172
rect -160 138 -148 172
rect -206 132 -148 138
rect -88 172 -30 178
rect -88 138 -76 172
rect -42 138 -30 172
rect -88 132 -30 138
rect 30 172 88 178
rect 30 138 42 172
rect 76 138 88 172
rect 30 132 88 138
rect 148 172 206 178
rect 148 138 160 172
rect 194 138 206 172
rect 148 132 206 138
rect 266 172 324 178
rect 266 138 278 172
rect 312 138 324 172
rect 266 132 324 138
rect 384 172 442 178
rect 384 138 396 172
rect 430 138 442 172
rect 384 132 442 138
rect 502 172 560 178
rect 502 138 514 172
rect 548 138 560 172
rect 502 132 560 138
rect -613 88 -567 100
rect -613 -88 -607 88
rect -573 -88 -567 88
rect -613 -100 -567 -88
rect -495 88 -449 100
rect -495 -88 -489 88
rect -455 -88 -449 88
rect -495 -100 -449 -88
rect -377 88 -331 100
rect -377 -88 -371 88
rect -337 -88 -331 88
rect -377 -100 -331 -88
rect -259 88 -213 100
rect -259 -88 -253 88
rect -219 -88 -213 88
rect -259 -100 -213 -88
rect -141 88 -95 100
rect -141 -88 -135 88
rect -101 -88 -95 88
rect -141 -100 -95 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 95 88 141 100
rect 95 -88 101 88
rect 135 -88 141 88
rect 95 -100 141 -88
rect 213 88 259 100
rect 213 -88 219 88
rect 253 -88 259 88
rect 213 -100 259 -88
rect 331 88 377 100
rect 331 -88 337 88
rect 371 -88 377 88
rect 331 -100 377 -88
rect 449 88 495 100
rect 449 -88 455 88
rect 489 -88 495 88
rect 449 -100 495 -88
rect 567 88 613 100
rect 567 -88 573 88
rect 607 -88 613 88
rect 567 -100 613 -88
rect -560 -138 -502 -132
rect -560 -172 -548 -138
rect -514 -172 -502 -138
rect -560 -178 -502 -172
rect -442 -138 -384 -132
rect -442 -172 -430 -138
rect -396 -172 -384 -138
rect -442 -178 -384 -172
rect -324 -138 -266 -132
rect -324 -172 -312 -138
rect -278 -172 -266 -138
rect -324 -178 -266 -172
rect -206 -138 -148 -132
rect -206 -172 -194 -138
rect -160 -172 -148 -138
rect -206 -178 -148 -172
rect -88 -138 -30 -132
rect -88 -172 -76 -138
rect -42 -172 -30 -138
rect -88 -178 -30 -172
rect 30 -138 88 -132
rect 30 -172 42 -138
rect 76 -172 88 -138
rect 30 -178 88 -172
rect 148 -138 206 -132
rect 148 -172 160 -138
rect 194 -172 206 -138
rect 148 -178 206 -172
rect 266 -138 324 -132
rect 266 -172 278 -138
rect 312 -172 324 -138
rect 266 -178 324 -172
rect 384 -138 442 -132
rect 384 -172 396 -138
rect 430 -172 442 -138
rect 384 -178 442 -172
rect 502 -138 560 -132
rect 502 -172 514 -138
rect 548 -172 560 -138
rect 502 -178 560 -172
rect -560 -246 -502 -240
rect -560 -280 -548 -246
rect -514 -280 -502 -246
rect -560 -286 -502 -280
rect -442 -246 -384 -240
rect -442 -280 -430 -246
rect -396 -280 -384 -246
rect -442 -286 -384 -280
rect -324 -246 -266 -240
rect -324 -280 -312 -246
rect -278 -280 -266 -246
rect -324 -286 -266 -280
rect -206 -246 -148 -240
rect -206 -280 -194 -246
rect -160 -280 -148 -246
rect -206 -286 -148 -280
rect -88 -246 -30 -240
rect -88 -280 -76 -246
rect -42 -280 -30 -246
rect -88 -286 -30 -280
rect 30 -246 88 -240
rect 30 -280 42 -246
rect 76 -280 88 -246
rect 30 -286 88 -280
rect 148 -246 206 -240
rect 148 -280 160 -246
rect 194 -280 206 -246
rect 148 -286 206 -280
rect 266 -246 324 -240
rect 266 -280 278 -246
rect 312 -280 324 -246
rect 266 -286 324 -280
rect 384 -246 442 -240
rect 384 -280 396 -246
rect 430 -280 442 -246
rect 384 -286 442 -280
rect 502 -246 560 -240
rect 502 -280 514 -246
rect 548 -280 560 -246
rect 502 -286 560 -280
rect -613 -330 -567 -318
rect -613 -506 -607 -330
rect -573 -506 -567 -330
rect -613 -518 -567 -506
rect -495 -330 -449 -318
rect -495 -506 -489 -330
rect -455 -506 -449 -330
rect -495 -518 -449 -506
rect -377 -330 -331 -318
rect -377 -506 -371 -330
rect -337 -506 -331 -330
rect -377 -518 -331 -506
rect -259 -330 -213 -318
rect -259 -506 -253 -330
rect -219 -506 -213 -330
rect -259 -518 -213 -506
rect -141 -330 -95 -318
rect -141 -506 -135 -330
rect -101 -506 -95 -330
rect -141 -518 -95 -506
rect -23 -330 23 -318
rect -23 -506 -17 -330
rect 17 -506 23 -330
rect -23 -518 23 -506
rect 95 -330 141 -318
rect 95 -506 101 -330
rect 135 -506 141 -330
rect 95 -518 141 -506
rect 213 -330 259 -318
rect 213 -506 219 -330
rect 253 -506 259 -330
rect 213 -518 259 -506
rect 331 -330 377 -318
rect 331 -506 337 -330
rect 371 -506 377 -330
rect 331 -518 377 -506
rect 449 -330 495 -318
rect 449 -506 455 -330
rect 489 -506 495 -330
rect 449 -518 495 -506
rect 567 -330 613 -318
rect 567 -506 573 -330
rect 607 -506 613 -330
rect 567 -518 613 -506
rect -560 -556 -502 -550
rect -560 -590 -548 -556
rect -514 -590 -502 -556
rect -560 -596 -502 -590
rect -442 -556 -384 -550
rect -442 -590 -430 -556
rect -396 -590 -384 -556
rect -442 -596 -384 -590
rect -324 -556 -266 -550
rect -324 -590 -312 -556
rect -278 -590 -266 -556
rect -324 -596 -266 -590
rect -206 -556 -148 -550
rect -206 -590 -194 -556
rect -160 -590 -148 -556
rect -206 -596 -148 -590
rect -88 -556 -30 -550
rect -88 -590 -76 -556
rect -42 -590 -30 -556
rect -88 -596 -30 -590
rect 30 -556 88 -550
rect 30 -590 42 -556
rect 76 -590 88 -556
rect 30 -596 88 -590
rect 148 -556 206 -550
rect 148 -590 160 -556
rect 194 -590 206 -556
rect 148 -596 206 -590
rect 266 -556 324 -550
rect 266 -590 278 -556
rect 312 -590 324 -556
rect 266 -596 324 -590
rect 384 -556 442 -550
rect 384 -590 396 -556
rect 430 -590 442 -556
rect 384 -596 442 -590
rect 502 -556 560 -550
rect 502 -590 514 -556
rect 548 -590 560 -556
rect 502 -596 560 -590
rect -560 -664 -502 -658
rect -560 -698 -548 -664
rect -514 -698 -502 -664
rect -560 -704 -502 -698
rect -442 -664 -384 -658
rect -442 -698 -430 -664
rect -396 -698 -384 -664
rect -442 -704 -384 -698
rect -324 -664 -266 -658
rect -324 -698 -312 -664
rect -278 -698 -266 -664
rect -324 -704 -266 -698
rect -206 -664 -148 -658
rect -206 -698 -194 -664
rect -160 -698 -148 -664
rect -206 -704 -148 -698
rect -88 -664 -30 -658
rect -88 -698 -76 -664
rect -42 -698 -30 -664
rect -88 -704 -30 -698
rect 30 -664 88 -658
rect 30 -698 42 -664
rect 76 -698 88 -664
rect 30 -704 88 -698
rect 148 -664 206 -658
rect 148 -698 160 -664
rect 194 -698 206 -664
rect 148 -704 206 -698
rect 266 -664 324 -658
rect 266 -698 278 -664
rect 312 -698 324 -664
rect 266 -704 324 -698
rect 384 -664 442 -658
rect 384 -698 396 -664
rect 430 -698 442 -664
rect 384 -704 442 -698
rect 502 -664 560 -658
rect 502 -698 514 -664
rect 548 -698 560 -664
rect 502 -704 560 -698
rect -613 -748 -567 -736
rect -613 -924 -607 -748
rect -573 -924 -567 -748
rect -613 -936 -567 -924
rect -495 -748 -449 -736
rect -495 -924 -489 -748
rect -455 -924 -449 -748
rect -495 -936 -449 -924
rect -377 -748 -331 -736
rect -377 -924 -371 -748
rect -337 -924 -331 -748
rect -377 -936 -331 -924
rect -259 -748 -213 -736
rect -259 -924 -253 -748
rect -219 -924 -213 -748
rect -259 -936 -213 -924
rect -141 -748 -95 -736
rect -141 -924 -135 -748
rect -101 -924 -95 -748
rect -141 -936 -95 -924
rect -23 -748 23 -736
rect -23 -924 -17 -748
rect 17 -924 23 -748
rect -23 -936 23 -924
rect 95 -748 141 -736
rect 95 -924 101 -748
rect 135 -924 141 -748
rect 95 -936 141 -924
rect 213 -748 259 -736
rect 213 -924 219 -748
rect 253 -924 259 -748
rect 213 -936 259 -924
rect 331 -748 377 -736
rect 331 -924 337 -748
rect 371 -924 377 -748
rect 331 -936 377 -924
rect 449 -748 495 -736
rect 449 -924 455 -748
rect 489 -924 495 -748
rect 449 -936 495 -924
rect 567 -748 613 -736
rect 567 -924 573 -748
rect 607 -924 613 -748
rect 567 -936 613 -924
rect -560 -974 -502 -968
rect -560 -1008 -548 -974
rect -514 -1008 -502 -974
rect -560 -1014 -502 -1008
rect -442 -974 -384 -968
rect -442 -1008 -430 -974
rect -396 -1008 -384 -974
rect -442 -1014 -384 -1008
rect -324 -974 -266 -968
rect -324 -1008 -312 -974
rect -278 -1008 -266 -974
rect -324 -1014 -266 -1008
rect -206 -974 -148 -968
rect -206 -1008 -194 -974
rect -160 -1008 -148 -974
rect -206 -1014 -148 -1008
rect -88 -974 -30 -968
rect -88 -1008 -76 -974
rect -42 -1008 -30 -974
rect -88 -1014 -30 -1008
rect 30 -974 88 -968
rect 30 -1008 42 -974
rect 76 -1008 88 -974
rect 30 -1014 88 -1008
rect 148 -974 206 -968
rect 148 -1008 160 -974
rect 194 -1008 206 -974
rect 148 -1014 206 -1008
rect 266 -974 324 -968
rect 266 -1008 278 -974
rect 312 -1008 324 -974
rect 266 -1014 324 -1008
rect 384 -974 442 -968
rect 384 -1008 396 -974
rect 430 -1008 442 -974
rect 384 -1014 442 -1008
rect 502 -974 560 -968
rect 502 -1008 514 -974
rect 548 -1008 560 -974
rect 502 -1014 560 -1008
<< properties >>
string FIXED_BBOX -704 -1093 704 1093
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.3 m 5 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
