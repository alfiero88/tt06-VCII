magic
tech sky130A
timestamp 1713266475
<< pwell >>
rect -656 -205 656 205
<< nmos >>
rect -558 -100 -358 100
rect -329 -100 -129 100
rect -100 -100 100 100
rect 129 -100 329 100
rect 358 -100 558 100
<< ndiff >>
rect -587 94 -558 100
rect -587 -94 -581 94
rect -564 -94 -558 94
rect -587 -100 -558 -94
rect -358 94 -329 100
rect -358 -94 -352 94
rect -335 -94 -329 94
rect -358 -100 -329 -94
rect -129 94 -100 100
rect -129 -94 -123 94
rect -106 -94 -100 94
rect -129 -100 -100 -94
rect 100 94 129 100
rect 100 -94 106 94
rect 123 -94 129 94
rect 100 -100 129 -94
rect 329 94 358 100
rect 329 -94 335 94
rect 352 -94 358 94
rect 329 -100 358 -94
rect 558 94 587 100
rect 558 -94 564 94
rect 581 -94 587 94
rect 558 -100 587 -94
<< ndiffc >>
rect -581 -94 -564 94
rect -352 -94 -335 94
rect -123 -94 -106 94
rect 106 -94 123 94
rect 335 -94 352 94
rect 564 -94 581 94
<< psubdiff >>
rect -638 170 -590 187
rect 590 170 638 187
rect -638 139 -621 170
rect 621 139 638 170
rect -638 -170 -621 -139
rect 621 -170 638 -139
rect -638 -187 -590 -170
rect 590 -187 638 -170
<< psubdiffcont >>
rect -590 170 590 187
rect -638 -139 -621 139
rect 621 -139 638 139
rect -590 -187 590 -170
<< poly >>
rect -558 136 -358 144
rect -558 119 -550 136
rect -366 119 -358 136
rect -558 100 -358 119
rect -329 136 -129 144
rect -329 119 -321 136
rect -137 119 -129 136
rect -329 100 -129 119
rect -100 136 100 144
rect -100 119 -92 136
rect 92 119 100 136
rect -100 100 100 119
rect 129 136 329 144
rect 129 119 137 136
rect 321 119 329 136
rect 129 100 329 119
rect 358 136 558 144
rect 358 119 366 136
rect 550 119 558 136
rect 358 100 558 119
rect -558 -119 -358 -100
rect -558 -136 -550 -119
rect -366 -136 -358 -119
rect -558 -144 -358 -136
rect -329 -119 -129 -100
rect -329 -136 -321 -119
rect -137 -136 -129 -119
rect -329 -144 -129 -136
rect -100 -119 100 -100
rect -100 -136 -92 -119
rect 92 -136 100 -119
rect -100 -144 100 -136
rect 129 -119 329 -100
rect 129 -136 137 -119
rect 321 -136 329 -119
rect 129 -144 329 -136
rect 358 -119 558 -100
rect 358 -136 366 -119
rect 550 -136 558 -119
rect 358 -144 558 -136
<< polycont >>
rect -550 119 -366 136
rect -321 119 -137 136
rect -92 119 92 136
rect 137 119 321 136
rect 366 119 550 136
rect -550 -136 -366 -119
rect -321 -136 -137 -119
rect -92 -136 92 -119
rect 137 -136 321 -119
rect 366 -136 550 -119
<< locali >>
rect -638 170 -590 187
rect 590 170 638 187
rect -638 139 -621 170
rect 621 139 638 170
rect -558 119 -550 136
rect -366 119 -358 136
rect -329 119 -321 136
rect -137 119 -129 136
rect -100 119 -92 136
rect 92 119 100 136
rect 129 119 137 136
rect 321 119 329 136
rect 358 119 366 136
rect 550 119 558 136
rect -581 94 -564 102
rect -581 -102 -564 -94
rect -352 94 -335 102
rect -352 -102 -335 -94
rect -123 94 -106 102
rect -123 -102 -106 -94
rect 106 94 123 102
rect 106 -102 123 -94
rect 335 94 352 102
rect 335 -102 352 -94
rect 564 94 581 102
rect 564 -102 581 -94
rect -558 -136 -550 -119
rect -366 -136 -358 -119
rect -329 -136 -321 -119
rect -137 -136 -129 -119
rect -100 -136 -92 -119
rect 92 -136 100 -119
rect 129 -136 137 -119
rect 321 -136 329 -119
rect 358 -136 366 -119
rect 550 -136 558 -119
rect -638 -170 -621 -139
rect 621 -170 638 -139
rect -638 -187 -590 -170
rect 590 -187 638 -170
<< viali >>
rect -550 119 -366 136
rect -321 119 -137 136
rect -92 119 92 136
rect 137 119 321 136
rect 366 119 550 136
rect -581 -94 -564 94
rect -352 -94 -335 94
rect -123 -94 -106 94
rect 106 -94 123 94
rect 335 -94 352 94
rect 564 -94 581 94
rect -550 -136 -366 -119
rect -321 -136 -137 -119
rect -92 -136 92 -119
rect 137 -136 321 -119
rect 366 -136 550 -119
<< metal1 >>
rect -556 136 -360 139
rect -556 119 -550 136
rect -366 119 -360 136
rect -556 116 -360 119
rect -327 136 -131 139
rect -327 119 -321 136
rect -137 119 -131 136
rect -327 116 -131 119
rect -98 136 98 139
rect -98 119 -92 136
rect 92 119 98 136
rect -98 116 98 119
rect 131 136 327 139
rect 131 119 137 136
rect 321 119 327 136
rect 131 116 327 119
rect 360 136 556 139
rect 360 119 366 136
rect 550 119 556 136
rect 360 116 556 119
rect -584 94 -561 100
rect -584 -94 -581 94
rect -564 -94 -561 94
rect -584 -100 -561 -94
rect -355 94 -332 100
rect -355 -94 -352 94
rect -335 -94 -332 94
rect -355 -100 -332 -94
rect -126 94 -103 100
rect -126 -94 -123 94
rect -106 -94 -103 94
rect -126 -100 -103 -94
rect 103 94 126 100
rect 103 -94 106 94
rect 123 -94 126 94
rect 103 -100 126 -94
rect 332 94 355 100
rect 332 -94 335 94
rect 352 -94 355 94
rect 332 -100 355 -94
rect 561 94 584 100
rect 561 -94 564 94
rect 581 -94 584 94
rect 561 -100 584 -94
rect -556 -119 -360 -116
rect -556 -136 -550 -119
rect -366 -136 -360 -119
rect -556 -139 -360 -136
rect -327 -119 -131 -116
rect -327 -136 -321 -119
rect -137 -136 -131 -119
rect -327 -139 -131 -136
rect -98 -119 98 -116
rect -98 -136 -92 -119
rect 92 -136 98 -119
rect -98 -139 98 -136
rect 131 -119 327 -116
rect 131 -136 137 -119
rect 321 -136 327 -119
rect 131 -139 327 -136
rect 360 -119 556 -116
rect 360 -136 366 -119
rect 550 -136 556 -119
rect 360 -139 556 -136
<< properties >>
string FIXED_BBOX -629 -178 629 178
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.0 l 2.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
