* NGSPICE file created from VCII-final.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_V5FT3Q a_n1116_n288# a_n1276_n374# a_n658_n288# a_n1174_n200#
+ a_716_n288# a_258_n288# a_200_n200# a_n716_n200# a_n258_n200# a_1116_n200# a_n200_n288#
+ a_658_n200#
X0 a_1116_n200# a_716_n288# a_658_n200# a_n1276_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=2
**devattr s=11600,458 d=23200,916
X1 a_200_n200# a_n200_n288# a_n258_n200# a_n1276_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
**devattr s=11600,458 d=11600,458
X2 a_n716_n200# a_n1116_n288# a_n1174_n200# a_n1276_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=2
**devattr s=23200,916 d=11600,458
X3 a_658_n200# a_258_n288# a_200_n200# a_n1276_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
**devattr s=11600,458 d=11600,458
X4 a_n258_n200# a_n658_n288# a_n716_n200# a_n1276_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
**devattr s=11600,458 d=11600,458
.ends

.subckt sky130_fd_pr__pfet_01v8_3HZ9VM w_n296_n719# a_n100_n597# a_100_n500# a_n158_n500#
X0 a_100_n500# a_n100_n597# a_n158_n500# w_n296_n719# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__nfet_01v8_EPHDNF a_1803_n100# a_n2421_n274# a_1345_n100# a_n29_n100#
+ a_887_n100# a_n1803_n188# a_429_n100# a_n1345_n188# a_1861_n188# a_n1861_n100# a_1403_n188#
+ a_n887_n188# a_2261_n100# a_n1403_n100# a_945_n188# a_n429_n188# a_n2319_n100# a_487_n188#
+ a_n2261_n188# a_n945_n100# a_29_n188# a_n487_n100#
X0 a_n1403_n100# a_n1803_n188# a_n1861_n100# a_n2421_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X1 a_887_n100# a_487_n188# a_429_n100# a_n2421_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X2 a_1345_n100# a_945_n188# a_887_n100# a_n2421_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X3 a_2261_n100# a_1861_n188# a_1803_n100# a_n2421_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=11600,516
X4 a_1803_n100# a_1403_n188# a_1345_n100# a_n2421_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X5 a_429_n100# a_29_n188# a_n29_n100# a_n2421_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X6 a_n1861_n100# a_n2261_n188# a_n2319_n100# a_n2421_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
**devattr s=11600,516 d=5800,258
X7 a_n487_n100# a_n887_n188# a_n945_n100# a_n2421_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X8 a_n945_n100# a_n1345_n188# a_n1403_n100# a_n2421_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
X9 a_n29_n100# a_n429_n188# a_n487_n100# a_n2421_n274# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
**devattr s=5800,258 d=5800,258
.ends

.subckt sky130_fd_pr__nfet_01v8_GSBCLJ a_n225_n909# a_n129_109# a_n369_21# a_n465_931#
+ a_447_109# a_399_21# a_n321_n909# a_n177_n87# a_n81_n997# a_n321_109# a_n509_109#
+ a_n33_n909# a_n509_n909# a_159_109# a_n369_n87# a_111_931# a_447_n909# a_351_109#
+ a_n33_109# a_n611_n1083# a_159_n909# a_303_n997# a_n225_109# a_303_931# a_n177_21#
+ a_255_n909# a_399_n87# a_n465_n997# a_207_21# a_351_n909# a_n417_n909# a_63_109#
+ a_n81_931# a_15_n87# a_15_21# a_111_n997# a_n417_109# a_n273_931# a_n129_n909# a_n273_n997#
+ a_255_109# a_207_n87# a_63_n909#
X0 a_n33_n909# a_n81_n997# a_n129_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X1 a_351_n909# a_303_n997# a_255_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X2 a_255_n909# a_207_n87# a_159_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X3 a_n33_109# a_n81_931# a_n129_109# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X4 a_n321_n909# a_n369_n87# a_n417_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X5 a_255_109# a_207_21# a_159_109# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X6 a_351_109# a_303_931# a_255_109# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X7 a_159_109# a_111_931# a_63_109# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X8 a_447_109# a_399_21# a_351_109# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=49600,1724
X9 a_n321_109# a_n369_21# a_n417_109# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X10 a_n225_109# a_n273_931# a_n321_109# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X11 a_159_n909# a_111_n997# a_63_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X12 a_n417_109# a_n465_931# a_n509_109# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
**devattr s=49600,1724 d=26400,866
X13 a_n129_109# a_n177_21# a_n225_109# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X14 a_n225_n909# a_n273_n997# a_n321_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X15 a_447_n909# a_399_n87# a_351_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=49600,1724
X16 a_63_n909# a_15_n87# a_n33_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X17 a_63_109# a_15_21# a_n33_109# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X18 a_n129_n909# a_n177_n87# a_n225_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
**devattr s=26400,866 d=26400,866
X19 a_n417_n909# a_n465_n997# a_n509_n909# a_n611_n1083# sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
**devattr s=49600,1724 d=26400,866
.ends

.subckt sky130_fd_pr__pfet_01v8_BDVWJN a_n129_n500# a_n465_n597# a_63_n500# a_n225_n500#
+ a_399_531# a_111_n597# a_n321_n500# a_n273_n597# a_15_531# a_n33_n500# a_n509_n500#
+ a_207_531# a_447_n500# a_n81_n597# a_n177_531# a_159_n500# a_255_n500# a_n369_531#
+ a_351_n500# a_n417_n500# a_303_n597# w_n647_n719#
X0 a_n33_n500# a_n81_n597# a_n129_n500# w_n647_n719# sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
**devattr s=33000,1066 d=33000,1066
X1 a_351_n500# a_303_n597# a_255_n500# w_n647_n719# sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
**devattr s=33000,1066 d=33000,1066
X2 a_255_n500# a_207_531# a_159_n500# w_n647_n719# sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
**devattr s=33000,1066 d=33000,1066
X3 a_n321_n500# a_n369_531# a_n417_n500# w_n647_n719# sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
**devattr s=33000,1066 d=33000,1066
X4 a_159_n500# a_111_n597# a_63_n500# w_n647_n719# sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
**devattr s=33000,1066 d=33000,1066
X5 a_n225_n500# a_n273_n597# a_n321_n500# w_n647_n719# sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
**devattr s=33000,1066 d=33000,1066
X6 a_447_n500# a_399_531# a_351_n500# w_n647_n719# sky130_fd_pr__pfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
**devattr s=33000,1066 d=62000,2124
X7 a_63_n500# a_15_531# a_n33_n500# w_n647_n719# sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
**devattr s=33000,1066 d=33000,1066
X8 a_n129_n500# a_n177_531# a_n225_n500# w_n647_n719# sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
**devattr s=33000,1066 d=33000,1066
X9 a_n417_n500# a_n465_n597# a_n509_n500# w_n647_n719# sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
**devattr s=62000,2124 d=33000,1066
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_RF5GSL a_n35_784# a_n165_n1346# a_n35_n1216#
X0 a_n35_784# a_n35_n1216# a_n165_n1346# sky130_fd_pr__res_xhigh_po_0p35 l=8
.ends

.subckt sky130_fd_pr__res_high_po_0p35_FFK5MY a_n35_n1416# a_n35_984# a_n165_n1546#
X0 a_n35_984# a_n35_n1416# a_n165_n1546# sky130_fd_pr__res_high_po_0p35 l=10
.ends

.subckt sky130_fd_pr__nfet_01v8_FMJ72H a_26_648# a_n383_n518# a_n147_n936# a_262_230#
+ a_498_648# a_n210_230# a_n210_n188# a_n446_648# a_n564_n188# a_207_n100# a_325_736#
+ a_n92_n606# a_380_n606# a_n446_n606# a_n29_318# a_n29_n100# a_443_n518# a_207_318#
+ a_207_n936# a_144_648# a_n265_n518# a_89_736# a_n210_n1024# a_n92_n1024# a_n92_n188#
+ a_n619_n518# a_n29_n936# a_n265_736# a_380_n188# a_n446_n188# a_n501_736# a_89_n100#
+ a_n147_318# a_262_n606# a_380_230# a_n328_n606# a_325_n518# a_144_n1024# a_n564_648#
+ a_n328_n1024# a_n147_n518# a_89_n936# a_n328_230# a_443_736# a_262_n188# a_n328_n188#
+ a_325_318# a_n92_230# a_262_648# a_n501_n100# a_n210_648# a_144_n606# a_498_n606#
+ a_207_n518# a_262_n1024# a_n446_n1024# a_n383_736# a_89_318# a_n501_n936# a_n29_n518#
+ a_n265_318# a_561_n100# a_n619_736# a_n501_318# a_144_n188# a_26_230# a_n383_n100#
+ a_498_n188# a_498_230# a_561_n936# a_n446_230# a_561_736# a_380_n1024# a_89_n518#
+ a_n564_n1024# a_n383_n936# a_26_n606# a_443_318# a_380_648# a_443_n100# a_144_230#
+ a_n265_n100# a_n328_648# a_n721_n1110# a_498_n1024# a_26_n188# a_n29_736# a_443_n936#
+ a_n619_n100# a_207_736# a_n383_318# a_n265_n936# a_n92_648# a_n501_n518# a_26_n1024#
+ a_n619_n936# a_n619_318# a_325_n100# a_n564_230# a_n147_n100# a_n210_n606# a_n147_736#
+ a_n564_n606# a_561_n518# a_561_318# a_325_n936#
X0 a_207_n100# a_144_n188# a_89_n100# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X1 a_89_n518# a_26_n606# a_n29_n518# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X2 a_207_n518# a_144_n606# a_89_n518# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X3 a_n29_n936# a_n92_n1024# a_n147_n936# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X4 a_n383_736# a_n446_648# a_n501_736# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X5 a_561_318# a_498_230# a_443_318# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=11600,516
X6 a_n29_736# a_n92_648# a_n147_736# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X7 a_325_318# a_262_230# a_207_318# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X8 a_n501_n100# a_n564_n188# a_n619_n100# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
**devattr s=11600,516 d=5800,258
X9 a_n501_n518# a_n564_n606# a_n619_n518# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
**devattr s=11600,516 d=5800,258
X10 a_n147_n518# a_n210_n606# a_n265_n518# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X11 a_325_n936# a_262_n1024# a_207_n936# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X12 a_n265_736# a_n328_648# a_n383_736# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X13 a_561_n936# a_498_n1024# a_443_n936# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=11600,516
X14 a_89_736# a_26_648# a_n29_736# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X15 a_207_318# a_144_230# a_89_318# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X16 a_n383_n100# a_n446_n188# a_n501_n100# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X17 a_n265_n936# a_n328_n1024# a_n383_n936# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X18 a_n147_736# a_n210_648# a_n265_736# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X19 a_n29_n100# a_n92_n188# a_n147_n100# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X20 a_443_n518# a_380_n606# a_325_n518# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X21 a_n501_318# a_n564_230# a_n619_318# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
**devattr s=11600,516 d=5800,258
X22 a_443_736# a_380_648# a_325_736# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X23 a_n265_n100# a_n328_n188# a_n383_n100# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X24 a_n383_n518# a_n446_n606# a_n501_n518# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X25 a_89_n936# a_26_n1024# a_n29_n936# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X26 a_207_n936# a_144_n1024# a_89_n936# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X27 a_561_736# a_498_648# a_443_736# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=11600,516
X28 a_n383_318# a_n446_230# a_n501_318# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X29 a_89_n100# a_26_n188# a_n29_n100# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X30 a_n29_n518# a_n92_n606# a_n147_n518# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X31 a_325_736# a_262_648# a_207_736# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X32 a_n501_n936# a_n564_n1024# a_n619_n936# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
**devattr s=11600,516 d=5800,258
X33 a_n147_n936# a_n210_n1024# a_n265_n936# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X34 a_n29_318# a_n92_230# a_n147_318# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X35 a_n147_n100# a_n210_n188# a_n265_n100# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X36 a_443_n100# a_380_n188# a_325_n100# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X37 a_325_n518# a_262_n606# a_207_n518# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X38 a_n265_318# a_n328_230# a_n383_318# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X39 a_207_736# a_144_648# a_89_736# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X40 a_561_n100# a_498_n188# a_443_n100# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=11600,516
X41 a_n265_n518# a_n328_n606# a_n383_n518# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X42 a_561_n518# a_498_n606# a_443_n518# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=11600,516
X43 a_89_318# a_26_230# a_n29_318# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X44 a_443_n936# a_380_n1024# a_325_n936# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X45 a_n501_736# a_n564_648# a_n619_736# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
**devattr s=11600,516 d=5800,258
X46 a_325_n100# a_262_n188# a_207_n100# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X47 a_n147_318# a_n210_230# a_n265_318# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X48 a_443_318# a_380_230# a_325_318# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
X49 a_n383_n936# a_n446_n1024# a_n501_n936# a_n721_n1110# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
**devattr s=5800,258 d=5800,258
.ends

.subckt sky130_fd_pr__pfet_01v8_3H5TVM a_158_n197# a_n416_n100# w_n812_n319# a_n358_n197#
+ a_358_n100# a_416_n197# a_n100_n197# a_100_n100# a_n674_n100# a_n158_n100# a_n616_n197#
+ a_616_n100#
X0 a_n158_n100# a_n358_n197# a_n416_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X1 a_100_n100# a_n100_n197# a_n158_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X2 a_616_n100# a_416_n197# a_358_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=11600,516
X3 a_358_n100# a_158_n197# a_100_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
**devattr s=5800,258 d=5800,258
X4 a_n416_n100# a_n616_n197# a_n674_n100# w_n812_n319# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
**devattr s=11600,516 d=5800,258
.ends

.subckt sky130_fd_pr__nfet_01v8_SMX62R a_n1209_n200# a_262_n288# a_n328_n288# a_1033_n200#
+ a_n501_n200# a_n855_n200# a_616_n288# a_561_n200# a_144_n288# a_n383_n200# a_498_n288#
+ a_915_n200# a_n1154_n288# a_n737_n200# a_443_n200# a_n1311_n374# a_797_n200# a_n265_n200#
+ a_n800_n288# a_n1036_n288# a_n619_n200# a_26_n288# a_325_n200# a_n682_n288# a_679_n200#
+ a_n147_n200# a_970_n288# a_n1091_n200# a_207_n200# a_n210_n288# a_n564_n288# a_852_n288#
+ a_n918_n288# a_n29_n200# a_380_n288# a_n92_n288# a_89_n200# a_n446_n288# a_1151_n200#
+ a_734_n288# a_n973_n200# a_1088_n288#
X0 a_n29_n200# a_n92_n288# a_n147_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X1 a_915_n200# a_852_n288# a_797_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X2 a_n619_n200# a_n682_n288# a_n737_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X3 a_n855_n200# a_n918_n288# a_n973_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X4 a_325_n200# a_262_n288# a_207_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X5 a_561_n200# a_498_n288# a_443_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X6 a_n265_n200# a_n328_n288# a_n383_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X7 a_1151_n200# a_1088_n288# a_1033_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=23200,916
X8 a_797_n200# a_734_n288# a_679_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X9 a_89_n200# a_26_n288# a_n29_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X10 a_207_n200# a_144_n288# a_89_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X11 a_n1091_n200# a_n1154_n288# a_n1209_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.3
**devattr s=23200,916 d=11600,458
X12 a_n501_n200# a_n564_n288# a_n619_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X13 a_n147_n200# a_n210_n288# a_n265_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X14 a_679_n200# a_616_n288# a_561_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X15 a_1033_n200# a_970_n288# a_915_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X16 a_n737_n200# a_n800_n288# a_n855_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X17 a_n973_n200# a_n1036_n288# a_n1091_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X18 a_443_n200# a_380_n288# a_325_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
X19 a_n383_n200# a_n446_n288# a_n501_n200# a_n1311_n374# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.3
**devattr s=11600,458 d=11600,458
.ends

.subckt sky130_fd_pr__pfet_01v8_P7N2DR a_2551_n250# a_n2351_486# a_n1061_1958# a_1319_1861#
+ a_2293_n986# a_2351_n1083# a_n1777_n347# a_n1777_n2555# a_n1835_486# a_n1835_n986#
+ a_29_n347# a_n1061_n1722# a_2351_n2555# a_n2351_n2458# a_1835_n1083# a_n2293_1861#
+ a_1261_n1722# a_1061_1861# a_2551_n2458# a_1777_n250# a_n2609_n250# a_1835_n2555#
+ a_n1835_n2458# a_n803_486# a_n1319_486# a_n2551_389# a_745_1958# a_n745_n347# a_1003_1222#
+ a_1835_1125# a_n229_n1083# a_n803_n986# a_n2035_n1819# a_n2609_n1722# a_1519_n986#
+ a_n2351_n250# a_2293_486# a_n229_n2555# a_1061_n1083# a_1777_486# a_n2035_389# a_n229_1125#
+ a_2551_1958# a_n1519_n1819# a_n2093_n986# a_1261_486# a_29_389# a_n1003_389# a_n1519_389#
+ a_n1003_1125# a_n1519_1861# a_1061_n2555# a_n1061_n2458# a_287_1125# a_803_n347#
+ a_n2035_n347# a_1261_n986# a_229_n250# a_1261_n2458# a_n2551_n1083# a_n1577_n250#
+ a_1777_1958# a_n487_1861# a_n2609_1958# a_745_486# a_2093_1125# a_n1261_1861# a_2035_n250#
+ a_545_n1819# a_2035_n1722# a_n2551_n2555# a_n487_n1819# a_29_n1819# a_n1319_n1722#
+ a_n29_1222# a_n2609_n2458# a_1519_n1722# a_n1319_n986# a_487_1222# a_n2351_1958#
+ a_229_486# a_545_1861# a_n545_n250# a_487_n1722# a_1835_n347# a_287_389# a_n287_n986#
+ a_2293_1222# a_n1061_n986# a_n2093_486# a_229_1958# a_2351_1861# a_n1261_n1083#
+ a_n229_n347# a_n1835_1222# a_n287_n1722# a_1319_n1083# a_n1061_486# a_n1577_486#
+ a_1319_1125# a_n1577_1958# a_n1003_n347# a_n1261_n2555# a_2035_n2458# a_1319_n2555#
+ a_287_n347# a_2035_1958# a_n1319_n2458# a_287_n1083# a_n2293_1125# a_n2293_389#
+ a_1519_n2458# a_n545_486# a_1061_1125# a_1577_1861# a_745_n986# a_1003_n250# a_n1777_389#
+ a_287_n2555# a_2093_n347# a_n1261_389# a_n803_1222# a_n545_1958# a_487_n2458# a_1519_1222#
+ a_2551_n986# a_2093_n1819# a_n2093_1222# a_n287_n2458# a_n745_389# a_1577_n1819#
+ a_n2551_1861# a_n1003_n1819# a_n745_n1819# a_803_n1819# a_1261_1222# a_n1519_1125#
+ a_n2035_n1083# a_1777_n986# a_n2609_n986# a_n1519_n1083# a_1319_n347# a_n229_389#
+ a_n2035_n2555# a_487_486# a_n487_1125# a_745_n1722# a_1003_1958# a_n1261_1125# a_n1777_1861#
+ a_n1519_n2555# a_n29_n250# a_n1319_1222# a_n2293_n347# a_29_1861# a_n2351_n986#
+ a_n545_n1722# a_487_n250# a_1061_n347# a_n29_486# a_1003_n1722# a_n287_1222# a_545_1125#
+ a_545_n1083# a_n1061_1222# a_29_n1083# a_n487_n1083# a_2293_n250# a_229_n986# a_n2293_n1819#
+ a_n745_1861# a_n1835_n250# a_2351_389# a_545_n2555# a_n1577_n986# a_2351_1125# a_n487_n2555#
+ a_29_n2555# a_1835_389# a_n1777_n1819# a_2035_n986# a_745_n2458# a_n1519_n347# a_2351_n1819#
+ a_n29_1958# a_745_1222# a_n287_486# a_n545_n2458# a_1319_389# a_487_1958# a_803_1861#
+ a_n2035_1861# a_1835_n1819# a_n803_n250# a_n487_n347# a_1577_1125# a_n545_n986#
+ a_n2093_n1722# a_1003_n2458# a_803_389# a_1519_n250# a_n1261_n347# a_2293_n1722#
+ a_2551_1222# a_n1577_n1722# a_n2093_n250# a_2293_1958# a_n487_389# a_n1835_1958#
+ a_n229_n1819# a_n29_n1722# a_1777_n1722# a_1261_n250# a_545_n347# a_n2609_486# a_n2551_1125#
+ a_1061_n1819# a_1777_1222# a_2093_n1083# a_n2609_1222# a_n803_n1722# a_1835_1861#
+ a_229_n1722# a_2351_n347# a_1003_n986# a_1577_n1083# a_n803_1958# a_2093_n2555#
+ a_n2093_n2458# a_803_n1083# a_n745_n1083# a_n1003_n1083# a_n229_1861# a_n1319_n250#
+ a_2551_486# a_1519_1958# w_n2747_n2677# a_n2551_n1819# a_2293_n2458# a_n2351_1222#
+ a_n1777_1125# a_1577_n2555# a_n1577_n2458# a_n2093_1958# a_n1003_1861# a_n1003_n2555#
+ a_n745_n2555# a_803_n2555# a_29_1125# a_287_1861# a_n29_n2458# a_1777_n2458# a_n287_n250#
+ a_1577_n347# a_n1061_n250# a_2035_486# a_229_1222# a_1261_1958# a_1519_486# a_1003_486#
+ a_2093_389# a_2093_1861# a_n803_n2458# a_n1577_1222# a_1577_389# a_n745_1125# a_229_n2458#
+ a_1061_389# a_n2351_n1722# a_2035_1222# a_2551_n1722# a_n29_n986# a_n1261_n1819#
+ a_n1835_n1722# a_n2551_n347# a_n1319_1958# a_1319_n1819# a_n2293_n1083# a_745_n250#
+ a_487_n986# a_n545_1222# a_803_1125# a_n2035_1125# a_287_n1819# a_n2293_n2555# a_n1777_n1083#
+ a_545_389# a_n287_1958#
X0 a_229_n1722# a_29_n1819# a_n29_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X1 a_n545_n1722# a_n745_n1819# a_n803_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X2 a_n1319_n986# a_n1519_n1083# a_n1577_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X3 a_229_n2458# a_29_n2555# a_n29_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X4 a_n545_n2458# a_n745_n2555# a_n803_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X5 a_n545_n986# a_n745_n1083# a_n803_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X6 a_2293_n986# a_2093_n1083# a_2035_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X7 a_n1577_1958# a_n1777_1861# a_n1835_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X8 a_n1061_n250# a_n1261_n347# a_n1319_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X9 a_1519_1958# a_1319_1861# a_1261_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X10 a_n287_n986# a_n487_n1083# a_n545_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X11 a_n2351_486# a_n2551_389# a_n2609_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=1
**devattr s=29000,1116 d=14500,558
X12 a_n803_n986# a_n1003_n1083# a_n1061_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X13 a_1003_n250# a_803_n347# a_745_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X14 a_n1061_1958# a_n1261_1861# a_n1319_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X15 a_n1577_1222# a_n1777_1125# a_n1835_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X16 a_1519_1222# a_1319_1125# a_1261_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X17 a_745_n250# a_545_n347# a_487_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X18 a_487_n250# a_287_n347# a_229_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X19 a_1003_1958# a_803_1861# a_745_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X20 a_1777_486# a_1577_389# a_1519_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X21 a_n1061_1222# a_n1261_1125# a_n1319_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X22 a_745_1958# a_545_1861# a_487_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X23 a_2293_486# a_2093_389# a_2035_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X24 a_487_1958# a_287_1861# a_229_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X25 a_1003_1222# a_803_1125# a_745_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X26 a_745_1222# a_545_1125# a_487_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X27 a_n2351_n1722# a_n2551_n1819# a_n2609_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=1
**devattr s=29000,1116 d=14500,558
X28 a_n2351_n2458# a_n2551_n2555# a_n2609_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=1
**devattr s=29000,1116 d=14500,558
X29 a_1003_n1722# a_803_n1819# a_745_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X30 a_487_1222# a_287_1125# a_229_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X31 a_1003_n2458# a_803_n2555# a_745_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X32 a_2035_n250# a_1835_n347# a_1777_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X33 a_1003_486# a_803_389# a_745_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X34 a_1777_n250# a_1577_n347# a_1519_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X35 a_n1577_n986# a_n1777_n1083# a_n1835_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X36 a_n1061_n1722# a_n1261_n1819# a_n1319_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X37 a_1519_n986# a_1319_n1083# a_1261_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X38 a_2035_1958# a_1835_1861# a_1777_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X39 a_n1577_486# a_n1777_389# a_n1835_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X40 a_n1061_n2458# a_n1261_n2555# a_n1319_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X41 a_1777_1958# a_1577_1861# a_1519_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X42 a_n2093_486# a_n2293_389# a_n2351_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X43 a_1261_n250# a_1061_n347# a_1003_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X44 a_n803_n1722# a_n1003_n1819# a_n1061_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X45 a_n803_n2458# a_n1003_n2555# a_n1061_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X46 a_n1061_n986# a_n1261_n1083# a_n1319_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X47 a_2035_1222# a_1835_1125# a_1777_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X48 a_n1835_n250# a_n2035_n347# a_n2093_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X49 a_1777_1222# a_1577_1125# a_1519_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X50 a_1261_1958# a_1061_1861# a_1003_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X51 a_1003_n986# a_803_n1083# a_745_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X52 a_745_n986# a_545_n1083# a_487_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X53 a_n1835_1958# a_n2035_1861# a_n2093_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X54 a_487_n986# a_287_n1083# a_229_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X55 a_1261_1222# a_1061_1125# a_1003_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X56 a_n1835_1222# a_n2035_1125# a_n2093_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X57 a_n803_486# a_n1003_389# a_n1061_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X58 a_745_486# a_545_389# a_487_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X59 a_n29_486# a_n229_389# a_n287_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X60 a_2035_n986# a_1835_n1083# a_1777_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X61 a_1777_n1722# a_1577_n1819# a_1519_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X62 a_1777_n986# a_1577_n1083# a_1519_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X63 a_1777_n2458# a_1577_n2555# a_1519_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X64 a_n2351_n250# a_n2551_n347# a_n2609_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=1
**devattr s=29000,1116 d=14500,558
X65 a_1519_n1722# a_1319_n1819# a_1261_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X66 a_1519_n2458# a_1319_n2555# a_1261_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X67 a_1261_n986# a_1061_n1083# a_1003_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X68 a_229_486# a_29_389# a_n29_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X69 a_n2093_n250# a_n2293_n347# a_n2351_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X70 a_229_n250# a_29_n347# a_n29_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X71 a_n1835_n986# a_n2035_n1083# a_n2093_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X72 a_n29_n250# a_n229_n347# a_n287_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X73 a_n2351_1958# a_n2551_1861# a_n2609_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=1
**devattr s=29000,1116 d=14500,558
X74 a_n2093_1958# a_n2293_1861# a_n2351_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X75 a_229_1958# a_29_1861# a_n29_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X76 a_n29_1958# a_n229_1861# a_n287_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X77 a_n2351_1222# a_n2551_1125# a_n2609_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=1
**devattr s=29000,1116 d=14500,558
X78 a_487_n1722# a_287_n1819# a_229_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X79 a_487_n2458# a_287_n2555# a_229_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X80 a_1519_486# a_1319_389# a_1261_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X81 a_2293_n1722# a_2093_n1819# a_2035_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X82 a_n2093_1222# a_n2293_1125# a_n2351_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X83 a_2293_n2458# a_2093_n2555# a_2035_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X84 a_229_1222# a_29_1125# a_n29_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X85 a_n29_1222# a_n229_1125# a_n287_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X86 a_487_486# a_287_389# a_229_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X87 a_n287_n1722# a_n487_n1819# a_n545_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X88 a_n287_n2458# a_n487_n2555# a_n545_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X89 a_n545_486# a_n745_389# a_n803_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X90 a_n1319_486# a_n1519_389# a_n1577_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X91 a_n29_n1722# a_n229_n1819# a_n287_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X92 a_n1577_n1722# a_n1777_n1819# a_n1835_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X93 a_2551_n250# a_2351_n347# a_2293_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=29000,1116
X94 a_n1319_n250# a_n1519_n347# a_n1577_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X95 a_n29_n2458# a_n229_n2555# a_n287_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X96 a_n1577_n2458# a_n1777_n2555# a_n1835_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X97 a_n1835_486# a_n2035_389# a_n2093_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X98 a_n2351_n986# a_n2551_n1083# a_n2609_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=1
**devattr s=29000,1116 d=14500,558
X99 a_2293_n250# a_2093_n347# a_2035_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X100 a_n545_n250# a_n745_n347# a_n803_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X101 a_2035_n1722# a_1835_n1819# a_1777_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X102 a_2035_n2458# a_1835_n2555# a_1777_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X103 a_n2093_n986# a_n2293_n1083# a_n2351_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X104 a_n287_n250# a_n487_n347# a_n545_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X105 a_n1319_n1722# a_n1519_n1819# a_n1577_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X106 a_2551_1958# a_2351_1861# a_2293_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=29000,1116
X107 a_n1319_n2458# a_n1519_n2555# a_n1577_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X108 a_229_n986# a_29_n1083# a_n29_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X109 a_n803_n250# a_n1003_n347# a_n1061_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X110 a_n1319_1958# a_n1519_1861# a_n1577_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X111 a_n29_n986# a_n229_n1083# a_n287_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X112 a_1261_486# a_1061_389# a_1003_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X113 a_n545_1958# a_n745_1861# a_n803_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X114 a_2293_1958# a_2093_1861# a_2035_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X115 a_n287_1958# a_n487_1861# a_n545_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X116 a_n1319_1222# a_n1519_1125# a_n1577_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X117 a_2551_1222# a_2351_1125# a_2293_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=29000,1116
X118 a_n803_1958# a_n1003_1861# a_n1061_1958# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X119 a_n545_1222# a_n745_1125# a_n803_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X120 a_2293_1222# a_2093_1125# a_2035_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X121 a_n287_1222# a_n487_1125# a_n545_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X122 a_n2093_n1722# a_n2293_n1819# a_n2351_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X123 a_2035_486# a_1835_389# a_1777_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X124 a_n803_1222# a_n1003_1125# a_n1061_1222# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X125 a_n2093_n2458# a_n2293_n2555# a_n2351_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X126 a_745_n1722# a_545_n1819# a_487_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X127 a_745_n2458# a_545_n2555# a_487_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X128 a_2551_n1722# a_2351_n1819# a_2293_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=29000,1116
X129 a_2551_486# a_2351_389# a_2293_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=29000,1116
X130 a_2551_n2458# a_2351_n2555# a_2293_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=29000,1116
X131 a_n1061_486# a_n1261_389# a_n1319_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X132 a_n1835_n2458# a_n2035_n2555# a_n2093_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X133 a_n1835_n1722# a_n2035_n1819# a_n2093_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X134 a_n287_486# a_n487_389# a_n545_486# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X135 a_1261_n1722# a_1061_n1819# a_1003_n1722# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X136 a_1261_n2458# a_1061_n2555# a_1003_n2458# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X137 a_n1577_n250# a_n1777_n347# a_n1835_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X138 a_1519_n250# a_1319_n347# a_1261_n250# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=14500,558
X139 a_2551_n986# a_2351_n1083# a_2293_n986# w_n2747_n2677# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=1
**devattr s=14500,558 d=29000,1116
.ends

.subckt VCII-final vdd vss z y ref x
XXM12 G2 vss G2 vss G2 G2 z z vss z G2 vss sky130_fd_pr__nfet_01v8_V5FT3Q
XXM13 vdd m1_17538_2386# vdd m1_17538_2386# sky130_fd_pr__pfet_01v8_3HZ9VM
XXM14 m1_17538_2386# vss vss m1_17538_2386# m1_17538_2386# G2 vss G2 G2 m1_17538_2386#
+ G2 G2 vss vss G2 G2 vss G2 G2 m1_17538_2386# G2 vss sky130_fd_pr__nfet_01v8_EPHDNF
XXM15 vdd z G4 G4 z G4 z G4 G4 z z vdd z vdd G4 G4 z vdd vdd vss vdd G4 vdd G4 G4
+ z G4 G4 G4 vdd vdd z G4 G4 G4 G4 vdd G4 z G4 z G4 z sky130_fd_pr__nfet_01v8_GSBCLJ
XXM16 vdd m1_17538_2386# G4 vdd sky130_fd_pr__pfet_01v8_3HZ9VM
XXM17 vss x vss G4 x x vss x x G4 vss x vss x x G4 vss x G4 G4 x G4 sky130_fd_pr__pfet_01v8_BDVWJN
XXR1 m1_1128_7074# vss m1_1502_5068# sky130_fd_pr__res_xhigh_po_0p35_RF5GSL
XXR2 m1_1128_7074# vss vdd sky130_fd_pr__res_xhigh_po_0p35_RF5GSL
XXR3 m1_1872_7070# vss m1_1502_5068# sky130_fd_pr__res_xhigh_po_0p35_RF5GSL
XXR4 m1_2290_5064# m1_1872_7070# vss sky130_fd_pr__res_high_po_0p35_FFK5MY
XXR5 G2 m1_2684_7472# vss sky130_fd_pr__res_high_po_0p35_FFK5MY
XXM1 ref G1 G1 ref ref ref ref ref ref B1 G1 ref ref ref B1 B1 B1 B1 B1 ref B1 G1
+ ref ref ref G1 B1 B1 ref ref B1 G1 G1 ref ref ref G1 ref ref ref G1 G1 ref B1 ref
+ ref G1 ref ref B1 ref ref ref B1 ref ref G1 G1 B1 B1 B1 G1 G1 B1 ref ref G1 ref
+ ref G1 ref G1 ref G1 ref G1 ref B1 ref B1 ref B1 ref vss ref ref B1 B1 G1 B1 G1
+ B1 ref B1 ref G1 G1 G1 ref G1 ref G1 ref G1 G1 G1 sky130_fd_pr__nfet_01v8_FMJ72H
XXR6 m1_2290_5064# m1_2684_7472# vss sky130_fd_pr__res_high_po_0p35_FFK5MY
XXM2 y D1 D1 y y y y y y B1 D1 y y y B1 B1 B1 B1 B1 y B1 D1 y y y D1 B1 B1 y y B1
+ D1 D1 y y y D1 y y y D1 D1 y B1 y y D1 y y B1 y y y B1 y y D1 D1 B1 B1 B1 D1 D1
+ B1 y y D1 y y D1 y D1 y D1 y D1 y B1 y B1 y B1 y vss y y B1 B1 D1 B1 D1 B1 y B1
+ y D1 D1 D1 y D1 y D1 y D1 D1 D1 sky130_fd_pr__nfet_01v8_FMJ72H
XXM3 G1 vdd vdd G1 D1 G1 G1 vdd D1 D1 G1 vdd sky130_fd_pr__pfet_01v8_3H5TVM
XXM4 G1 G1 vdd G1 vdd G1 G1 G1 vdd vdd G1 G1 sky130_fd_pr__pfet_01v8_3H5TVM
XXM5 vss vss B1 vss vss G2 B1 G2 G2 vss G2 G2 B1 B1 G2 G2 B1 G2 G2 vss G2 B1 sky130_fd_pr__nfet_01v8_EPHDNF
XXM6 G2 vss vss G2 G2 G2 vss G2 G2 G2 G2 G2 vss vss G2 G2 vss G2 G2 G2 G2 vss sky130_fd_pr__nfet_01v8_EPHDNF
XXM7 y D1 D1 m1_7898_5534# y m1_7898_5534# D1 m1_7898_5534# D1 m1_7898_5534# D1 y
+ D1 y y vss m1_7898_5534# y D1 D1 m1_7898_5534# D1 m1_7898_5534# D1 y m1_7898_5534#
+ D1 m1_7898_5534# y D1 D1 D1 D1 y D1 D1 m1_7898_5534# D1 y D1 y D1 sky130_fd_pr__nfet_01v8_SMX62R
XXM8 y vss vss y y G2 vss G2 G2 y G2 G2 vss vss G2 G2 vss G2 G2 y G2 vss sky130_fd_pr__nfet_01v8_EPHDNF
XXM9 vdd m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# vdd m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd vdd m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ vdd m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# vdd m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# vdd vdd vdd m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ vdd vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd vdd m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ vdd vdd m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534#
+ vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd vdd m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# vdd vdd vdd vdd m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ vdd m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd vdd m1_7898_5534# vdd
+ vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# vdd
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ vdd vdd vdd m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# vdd vdd vdd m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd vdd vdd m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd vdd m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# vdd vdd m1_7898_5534# m1_7898_5534# vdd vdd m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ vdd vdd vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# vdd vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# sky130_fd_pr__pfet_01v8_P7N2DR
XXM10 vdd x vdd m1_7898_5534# x m1_7898_5534# m1_7898_5534# m1_7898_5534# x x m1_7898_5534#
+ vdd m1_7898_5534# x m1_7898_5534# m1_7898_5534# x m1_7898_5534# vdd x vdd m1_7898_5534#
+ x x x m1_7898_5534# x m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# x m1_7898_5534#
+ vdd vdd x x m1_7898_5534# m1_7898_5534# x m1_7898_5534# m1_7898_5534# vdd m1_7898_5534#
+ vdd x m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# x x x m1_7898_5534# vdd x m1_7898_5534#
+ vdd x m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# vdd m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# x vdd vdd vdd x vdd x x m1_7898_5534# vdd vdd m1_7898_5534# m1_7898_5534#
+ x x vdd vdd x m1_7898_5534# m1_7898_5534# m1_7898_5534# x x m1_7898_5534# vdd vdd
+ m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# vdd
+ x m1_7898_5534# m1_7898_5534# m1_7898_5534# vdd vdd m1_7898_5534# m1_7898_5534#
+ x vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# x vdd vdd vdd vdd
+ m1_7898_5534# vdd x m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# x m1_7898_5534# m1_7898_5534# x vdd m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# vdd m1_7898_5534# x vdd m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ vdd x m1_7898_5534# m1_7898_5534# x vdd vdd m1_7898_5534# vdd vdd x m1_7898_5534#
+ m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# x x m1_7898_5534# m1_7898_5534# x
+ m1_7898_5534# m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# vdd x m1_7898_5534# m1_7898_5534# vdd x x vdd m1_7898_5534# vdd m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# x m1_7898_5534# m1_7898_5534# vdd vdd vdd m1_7898_5534#
+ vdd m1_7898_5534# x vdd vdd vdd x m1_7898_5534# x m1_7898_5534# vdd x x m1_7898_5534#
+ vdd m1_7898_5534# m1_7898_5534# x m1_7898_5534# vdd x m1_7898_5534# x m1_7898_5534#
+ vdd m1_7898_5534# x m1_7898_5534# vdd m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# x vdd vdd vdd m1_7898_5534# x x m1_7898_5534# m1_7898_5534# vdd vdd
+ m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ vdd x x m1_7898_5534# vdd vdd x x vdd vdd m1_7898_5534# m1_7898_5534# x vdd m1_7898_5534#
+ m1_7898_5534# x m1_7898_5534# x vdd vdd vdd m1_7898_5534# x m1_7898_5534# x m1_7898_5534#
+ m1_7898_5534# x vdd vdd m1_7898_5534# m1_7898_5534# m1_7898_5534# m1_7898_5534#
+ m1_7898_5534# m1_7898_5534# x sky130_fd_pr__pfet_01v8_P7N2DR
XXM11 x vss vss x x G2 vss G2 G2 x G2 G2 vss vss G2 G2 vss G2 G2 x G2 vss sky130_fd_pr__nfet_01v8_EPHDNF
.ends

